* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65u l = 0.15u m = 2 ad = 0.231p pd = 1.93u as = 0.462p ps = 3.86u nrd = 240.00 nrs = 120.00 mult = {2*mult}
xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65u l = 0.15u m = 2 ad = 0.495p pd = 3.9u as = 0.0p ps = 0.0u nrd = 120.0 nrs = 0.0 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65u l = 0.15u m = 4 ad = 0.231p pd = 1.93u as = 0.347p ps = 2.90u nrd = 240.00 nrs = 160.00 mult = {4*mult}
xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65u l = 0.15u m = 2 ad = 0.495p pd = 3.9u as = 0.0p ps = 0.0u nrd = 120.00 nrs = 0.0 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65u l = 0.18u m = 2 ad = 0.231p pd = 1.93u as = 0.462p ps = 3.86u nrd = 240.00 nrs = 120.00 mult = {2*mult}
xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65u l = 0.18u m = 2 ad = 0.495p pd = 3.9u as = 0.0p ps = 0.0u nrd = 120.00 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p18
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65u l = 0.18u m = 4 ad = 0.231p pd = 1.93u as = 0.347p ps = 2.90u nrd = 240.00 nrs = 160.00 mult = {4*mult}
xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65u l = 0.18u m = 2 ad = 0.495p pd = 3.9u as = 0.0p ps = 0.0u nrd = 120.00 nrs = 0.0 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p18
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65u l = 0.25u m = 2 ad = 0.231p pd = 1.93u as = 0.462p ps = 3.86u nrd = 240.00 nrs = 120.00 mult = {2*mult}
xsky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02 w = 1.65u l = 0.25u m = 2 ad = 0.495p pd = 3.9u as = 0.0p ps = 0.0u nrd = 120.00 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM02W1p65L0p25
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65u l = 0.25u m = 4 ad = 0.231p pd = 1.93u as = 0.347p ps = 2.90u nrd = 240.00 nrs = 160.00 mult = {4*mult}
xsky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04 w = 1.65u l = 0.25u m = 2 ad = 0.495p pd = 3.9u as = 0.0p ps = 0.0u nrd = 120.00 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM04W1p65L0p25
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.15u m = 2 ad = 0.421p pd = 3.29u as = 0.843p ps = 6.58u nrd = 133.33 nrs = 66.67 mult = {2*mult}
xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.15u m = 2 ad = 0.903p pd = 6.62u as = 0.0p ps = 0.0u nrd = 66.67 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.15u m = 4 ad = 0.421p pd = 3.29u as = 0.632p ps = 4.94u nrd = 133.33 nrs = 88.89 mult = {4*mult}
xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.15u m = 2 ad = 0.903p pd = 6.62u as = 0.0p ps = 0.0u nrd = 66.67 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.18u m = 2 ad = 0.421p pd = 3.29u as = 0.843p ps = 6.58u nrd = 133.33 nrs = 66.67 mult = {2*mult}
xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.18u m = 2 ad = 0.903p pd = 6.62u as = 0.0p ps = 0.0u nrd = 66.67 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p18
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.18u m = 4 ad = 0.421p pd = 3.29u as = 0.632p ps = 4.94u nrd = 133.33 nrs = 88.89 mult = {4*mult}
xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.18u m = 2 ad = 0.903p pd = 6.62u as = 0.0p ps = 0.0u nrd = 66.67 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p18
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.25u m = 2 ad = 0.421p pd = 3.29u as = 0.843p ps = 6.58u nrd = 133.33 nrs = 66.67 mult = {2*mult}
xsky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W3p00 l = 0.25u m = 2 ad = 0.903p pd = 6.62u as = 0.0p ps = 0.0u nrd = 66.67 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM02W3p00L0p25
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.25u m = 4 ad = 0.421p pd = 3.29u as = 0.632p ps = 4.94u nrd = 133.33 nrs = 88.89 mult = {4*mult}
xsky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W3p00 l = 0.25u m = 2 ad = 0.903p pd = 6.62u as = 0.0p ps = 0.0u nrd = 66.67 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM04W3p00L0p25
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.15u m = 2 ad = 0.707p pd = 5.33u as = 1.414p ps = 10.66u nrd = 80.00 nrs = 40.00 mult = {2*mult}
xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.15u m = 2 ad = 1.515p pd = 10.7u as = 0.0p ps = 0.0u nrd = 40.00 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.15u m = 4 ad = 0.707p pd = 5.33u as = 1.061p ps = 8.00u nrd = 80.00 nrs = 53.33 mult = {4*mult}
xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.15u m = 2 ad = 1.515p pd = 10.7u as = 0.0p ps = 0.0u nrd = 40.00 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.18u m = 2 ad = 0.707p pd = 5.33u as = 1.414p ps = 10.66u nrd = 80.00 nrs = 40.00 mult = {2*mult}
xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.18u m = 2 ad = 1.515p pd = 10.7u as = 0.0p ps = 0.0u nrd = 40.00 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p18
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.18u m = 4 ad = 0.707p pd = 5.33u as = 1.061p ps = 8.00u nrd = 80.00 nrs = 53.33 mult = {4*mult}
xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.18u m = 2 ad = 1.515p pd = 10.7u as = 0.0p ps = 0.0u nrd = 40.00 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p18
.subckt  sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.25u m = 2 ad = 0.707p pd = 5.33u as = 1.414p ps = 10.66u nrd = 80.00 nrs = 40.00 mult = {2*mult}
xsky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM02W5p00 l = 0.25u m = 2 ad = 1.515p pd = 10.7u as = 0.0p ps = 0.0u nrd = 40.00 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25
.subckt  sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25 d g s b
+ 
.param  mult = 1.0
xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25 d g s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.25u m = 4 ad = 0.707p pd = 5.33u as = 1.061p ps = 8.00u nrd = 80.00 nrs = 53.33 mult = {4*mult}
xsky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25_dummy b b s b sky130_fd_pr__rf_pfet_01v8_bM04W5p00 l = 0.25u m = 2 ad = 1.515p pd = 10.7u as = 0.0p ps = 0.0u nrd = 40.00 nrs = 0.00 mult = {2*mult}
.ends sky130_fd_pr__rf_pfet_01v8_bM04W5p00L0p25
.subckt  sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15 d g s b
+ 
+ 
.param  mult = 1.0
+ rg_sub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult)}
+ rg_dist_tnom = {(150.129*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult)}
+ tref = 30.0
xsky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15u w = {(2)*(1.68u)} ad = {(2)*(0.2352p)} as = {(2)*(0.445p)} pd = {(2)*(1.96u)} ps = {(2)*(3.89u)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265u sb = 0.265u sd = 0.28u m = 1 mult = {1*mult}
cpar_ds 1  3 c = {(0.41f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
cpar_gd 2  1 c = {(0.74f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
cpar_gs 2  3 c = {(0.119f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
rg 2  g r = {(rg_sub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}
rd 1  d r = {(154*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}
rs 3  s r = {(76*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}
.ends sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15 d g s b
+ 
+ 
.param  mult = 1.0
+ rg_stub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2)}
+ rg_dist_tnom = {(366.81*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2)}
+ tref = 30.0
xsky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15u w = {(2)*(5.00u)} ad = {(2)*(0.7p)} as = {(2)*(1.325p)} pd = {(2)*(5.28u)} ps = {(2)*(10.53u)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265u sb = 0.265u sd = 0.28u m = 1 mult = {1*mult}
cpar_ds 1  3 c = {(1.22f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2)}
cpar_gd 2  1 c = {(1.665f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2)}
cpar_gs 2  3 c = {(0.285f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2)}
rg 2  g r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}
rd 1  d r = {(50*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}
rs 3  s r = {(24*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}
.ends sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15 d g s b
+ 
+ 
.param  mult = 1.0
+ rg_stub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2)}
+ rg_dist_tnom = {(37.53*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2)}
+ tref = 30.0
xsky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15u w = {(2)*(0.84u)} ad = {(2)*(0.1176p)} as = {(2)*(0.223p)} pd = {(2)*(1.12u)} ps = {(2)*(2.21u)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265u sb = 0.265u sd = 0.28u m = 1 mult = {1*mult}
cpar_ds 1  3 c = {(0.17f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
cpar_gd 2  1 c = {(0.459f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
cpar_gs 2  3 c = {(0.257f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
rg 2  g r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}
rd 1  d r = {(306*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}
rs 3  s r = {(152.5*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}
.ends sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15 d g s b
+ 
+ 
.param  mult = 1.0
+ rg_stub_tnom = {(63.5*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult)}
+ rg_dist_tnom = {(75.061*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult)}
+ tref = 30.0
xsky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15u w = {(4)*(1.68u)} ad = {(4)*(0.2352p)} as = {(4)*(0.34p)} pd = {(4)*(1.96u)} ps = {(4)*(2.925u)} nrd = {(0)/(4)} nrs = {(0)/(4)} nf = 4 sa = 0.265u sb = 0.265u sd = 0.28u m = 1 mult = {1*mult}
cpar_ds 1  3 c = {(0.82f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
cpar_gd 2  1 c = {(0.984f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
cpar_gs 2  3 c = {(0.354f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
rg 2  g r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}
rd 1  d r = {(78*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}
rs 3  s r = {(50.6*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}
.ends sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15
.subckt  sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15 d g s b
+ 
+ 
.param  mult = 1.0
+ rg_stub_tnom = {(127*sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult)}
+ rg_dist_tnom = {(183.0*sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult)}
+ tref = 30.0
xsky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15 1 2 3 b sky130_fd_pr__pfet_01v8 l = 0.15u w = {(2)*(3.00u)} ad = {(2)*(0.42p)} as = {(2)*(0.795p)} pd = {(2)*(3.28u)} ps = {(2)*(6.53u)} nrd = {(0)/(2)} nrs = {(0)/(2)} nf = 2 sa = 0.265u sb = 0.265u sd = 0.28u m = 1 mult = {1*mult}
cpar_ds 1  3  c = {(0.7f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
cpar_gd 2  1  c = {(1.056f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
cpar_gs 2  3  c = {(0.232f*sky130_fd_pr__rf_pfet_01v8__aw_cap_mult)}
rg 2  g  r = {(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))}
rd 1  d  r = {(78*sky130_fd_pr__rf_pfet_01v8__aw_rd_mult)}
rs 3  s  r = {(38.5*sky130_fd_pr__rf_pfet_01v8__aw_rs_mult)}
.ends sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15
