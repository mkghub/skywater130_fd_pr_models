* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 18
.param
+ sky130_fd_pr__rf_nfet_01v8_b__toxe_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_b__overlap_mult = 0.9642
+ sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult = 9.9543e-1
+ sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult = 1.0204
+ sky130_fd_pr__rf_nfet_01v8_b__lint_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_b__wint_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_b__rshg_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_b__dlc_diff = -.61492e-9
+ sky130_fd_pr__rf_nfet_01v8_b__dwc_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_b__xgw_diff = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_0 = -0.019045
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_0 = 876.33
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_0 = 0.0076402
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_0 = 0.00078682
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_0 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_1 = -0.0024718
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_1 = 292.74
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_1 = 0.01684
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_1 = 0.00069507
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_1 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_2 = -0.011464
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_2 = 4008.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_2 = 0.034561
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_2 = -0.00018668
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_2 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_3 = 0.0031296
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_3 = -7677.3
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_3 = 0.0045864
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_3 = -0.0050888
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_3 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_4 = -0.019118
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_4 = -3226.1
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_4 = 0.020455
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_4 = -0.0033825
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_4 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_5 = -0.010928
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_5 = -3103.8
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_5 = 0.037245
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_5 = -0.00010837
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_6 = -0.0038131
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_6 = -0.010357
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_6 = -10521.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_6 = 0.0019487
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_7 = 0.017771
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_7 = -0.0036526
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_7 = -0.018633
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_7 = -3856.6
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_7 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM02__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__k2_diff_8 = 0.03546
+ sky130_fd_pr__rf_nfet_01v8_bM02__u0_diff_8 = -0.0023259
+ sky130_fd_pr__rf_nfet_01v8_bM02__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM02__vth0_diff_8 = -0.014738
+ sky130_fd_pr__rf_nfet_01v8_bM02__vsat_diff_8 = -749.49
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_0 = 0.0066076
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_0 = -0.00069668
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_0 = 0.0055162
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_0 = -9578.4
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_0 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_1 = 0.022438
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_1 = -0.0013475
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_1 = -0.017125
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_1 = -1947.1
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_1 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_2 = 0.0375
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_2 = -0.0010013
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_2 = -0.013525
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_2 = 3934.3
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_3 = -9286.3
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_3 = 0.0055484
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_3 = -0.005738
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_3 = -0.0050065
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_3 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_4 = -2375.7
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_4 = 0.023623
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_4 = -0.0067253
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_4 = -0.025509
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_4 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_5 = 14291.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_5 = 0.039092
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_5 = -0.0049774
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_5 = -0.018429
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_5 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_6 = -11321.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_6 = 0.0029951
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_6 = -0.0037175
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_6 = -0.011302
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_7 = -0.0055361
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_7 = -8608.4
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_7 = 0.021579
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_7 = -0.029895
*
* sky130_fd_pr__rf_nfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_bM04__vth0_diff_8 = -0.019214
+ sky130_fd_pr__rf_nfet_01v8_bM04__u0_diff_8 = -0.0040927
+ sky130_fd_pr__rf_nfet_01v8_bM04__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__vsat_diff_8 = 9127.9
+ sky130_fd_pr__rf_nfet_01v8_bM04__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_bM04__k2_diff_8 = 0.037329
.include "sky130_fd_pr_models/cells/sky130_fd_pr__rf_nfet_01v8_b.pm3.spice"
