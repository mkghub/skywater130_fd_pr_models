* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__res_generic_po__slope = 0.0
.param sky130_fd_pr__res_generic_po__tc1_slope = 1.0
.param sky130_fd_pr__res_generic_po__tc2_slope = 1.0
* statistics {
*   mismatch {
*     vary  sky130_fd_pr__res_generic_po__slope dist=gauss std=0.12
*   }
*   process {
*     vary  sky130_fd_pr__res_generic_po__tc1_slope dist=gauss std=0.125
*     vary  sky130_fd_pr__res_generic_po__tc2_slope dist=gauss std=0.125
*   }
* }
.subckt  sky130_fd_pr__res_generic_po r0 r1
+ 
.param  w = 1u l = 0u mult = 1 r = 0 tc1 = {tc1rsgpu*sky130_fd_pr__res_generic_po__tc1_slope} tc2 = {tc2rsgpu*sky130_fd_pr__res_generic_po__tc2_slope}
+ rp1_mm = {rp1*sky130_fd_pr__res_generic_po__slope/sqrt(2.0*l*w*mult+rp1/100000.0)}
+ r_tot = {(rp1+rp1_mm)*l/(w-1e6*(-tol_poly-poly_dw))+r}
sky130_fd_pr__res_generic_po r0 r1 sky130_fd_pr__res_generic_po__monte r = {r_tot} tc1r = {tc1} tc2r = {tc2}
.model sky130_fd_pr__res_generic_po__monte r tref = 30.0
.ends sky130_fd_pr__res_generic_po
