* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 18
.param
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42 = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42 = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42 = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult = 1.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_0 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_1 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_2 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_3 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_4 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_5 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_6 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_7 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_8 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_0 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_1 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_2 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_3 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_4 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_5 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_6 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_7 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_8 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"
