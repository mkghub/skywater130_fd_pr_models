* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 68
.param
+ sky130_fd_pr__pfet_01v8_hvt__toxe_mult = 1.0365
+ sky130_fd_pr__pfet_01v8_hvt__rshp_mult = 1.0
+ sky130_fd_pr__pfet_01v8_hvt__overlap_mult = 1.1614
+ sky130_fd_pr__pfet_01v8_hvt__lint_diff = -1.21275e-8
+ sky130_fd_pr__pfet_01v8_hvt__wint_diff = 2.252e-8
+ sky130_fd_pr__pfet_01v8_hvt__dlc_diff = -1.21275e-8
+ sky130_fd_pr__pfet_01v8_hvt__dwc_diff = 2.252e-8
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 000, W = 1.26u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0 = -0.34579
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_0 = 0.020851
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_0 = -0.0095877
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_0 = 1.1114e-19
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_0 = 0.00034006
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0 = -5725.7
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0 = 0.034024
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_0 = 8.2585e-11
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 001, W = 1.68u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1 = 0.2871
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_1 = 0.028366
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_1 = -2.2775e-19
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_1 = -0.015152
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_1 = 0.0013261
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1 = -29348.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1 = 0.032845
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_1 = 4.1588e-10
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 002, W = 1.0u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2 = -0.046804
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_2 = 0.10489
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_2 = -0.16129
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_2 = -0.03535
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_2 = 1.174e-18
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_2 = -0.0094251
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_2 = 0.0030692
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2 = -0.048378
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_2 = -2.1209e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 003, W = 1.0u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_3 = -1.424e-10
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3 = 0.12144
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_3 = 0.041944
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_3 = -0.049051
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_3 = -0.023404
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_3 = 7.0752e-19
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_3 = -0.010721
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_3 = 0.0017002
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3 = -0.02632
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 004, W = 1.0u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_4 = -1.2493e-10
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4 = 0.099998
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_4 = 0.0049331
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_4 = -0.0098663
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_4 = -0.034079
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_4 = 6.9913e-19
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_4 = -0.011492
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_4 = 0.0019259
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4 = -0.028711
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_4 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 005, W = 1.0u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_5 = -1.6364e-11
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5 = 0.21275
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_5 = 0.078419
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_5 = -0.079421
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_5 = -0.033475
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_5 = 6.9612e-19
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_5 = -0.012817
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_5 = 0.0026926
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5 = -0.028045
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 006, W = 1.0u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_6 = 3.4181e-10
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6 = 0.5689
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_6 = -0.027227
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_6 = -2.4777e-19
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_6 = -0.027088
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_6 = 0.00096443
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6 = -3467.4
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6 = 0.0069854
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 007, W = 1.0u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_7 = -0.0010034
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_7 = 3.6357e-19
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7 = 36008.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7 = -0.01276
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_7 = -4.1129e-10
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7 = -0.31412
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_7 = 0.03096
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_7 = -0.010589
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 008, W = 1.0u, L = 0.25u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_8 = -0.013407
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_8 = -0.00058228
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_8 = -8.5158e-19
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8 = -42889.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8 = -0.037881
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_8 = 6.5523e-10
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8 = 0.43597
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_8 = -0.011121
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 009, W = 1.0u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_9 = -0.033668
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_9 = -0.0036582
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_9 = -0.0012153
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_9 = 9.1948e-19
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9 = 140000.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9 = -0.026553
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_9 = -7.8144e-10
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9 = -1.4
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 010, W = 3.0u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_10 = 2.6144e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_10 = -0.020127
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_10 = -0.0030239
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_10 = 0.0093741
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10 = 0.064133
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_10 = 0.0007345
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10 = -0.013796
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_10 = -0.011062
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_10 = -4.6435e-11
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 011, W = 3.0u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_11 = -7.1725e-11
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_11 = 3.6998e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_11 = -0.032292
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_11 = 0.0034784
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_11 = -0.0077387
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11 = 0.10742
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_11 = 0.001108
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11 = -0.017098
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_11 = -0.012484
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 012, W = 3.0u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_12 = -0.00081443
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_12 = -8.5857e-12
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_12 = 6.4556e-20
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_12 = 0.013024
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_12 = -0.0043204
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_12 = 0.0044821
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12 = 1.097
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_12 = 0.00034554
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12 = -0.0090812
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 013, W = 3.0u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13 = 1.1856
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_13 = 0.000291
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13 = 0.0013183
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_13 = -0.0030908
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_13 = -8.0647e-12
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_13 = 7.1302e-20
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_13 = 0.0050583
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_13 = -0.0097395
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_13 = 0.0067576
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 014, W = 3.0u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14 = -24055.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14 = -0.045104
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_14 = 0.00083795
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14 = 0.044387
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_14 = -0.011007
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_14 = 1.2431e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_14 = 1.1518e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_14 = 0.0072954
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_14 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 015, W = 3.0u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15 = 10640.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15 = 0.35651
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_15 = 0.001258
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15 = 0.0073327
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_15 = -0.019393
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_15 = 1.795e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_15 = 1.4895e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_15 = -0.027125
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_15 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 016, W = 3.0u, L = 0.25u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16 = -2684.8
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16 = 0.4167
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_16 = 0.00094935
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16 = -0.033644
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_16 = -6.0646e-5
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_16 = 1.0769e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_16 = 2.9025e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_16 = -0.0094744
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 017, W = 3.0u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17 = -0.071718
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_17 = 0.00057944
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17 = 19087.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17 = -0.012025
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_17 = -0.0082116
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_17 = 6.4163e-11
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_17 = 1.0541e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_17 = -0.01648
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_17 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 018, W = 5.0u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_18 = 0.011929
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_18 = -0.015714
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18 = 0.051526
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_18 = 0.00092609
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18 = -0.013451
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_18 = -0.01165
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_18 = -5.9564e-11
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_18 = 3.3986e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_18 = -0.023431
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 019, W = 5.0u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_19 = -0.01949
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_19 = -0.0027099
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_19 = 0.0037748
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19 = 0.077586
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_19 = -6.633e-5
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19 = -0.0033747
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_19 = -0.0056173
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_19 = -2.0295e-12
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_19 = -1.1262e-20
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 020, W = 5.0u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_20 = -0.0016805
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_20 = -0.040992
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_20 = 0.04802
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20 = 0.017444
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_20 = -0.00019237
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20 = 0.0062824
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_20 = -0.0012963
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_20 = 3.6986e-11
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_20 = -8.1372e-20
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 021, W = 5.0u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_21 = -3.5987e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_21 = 0.01627
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_21 = -0.10035
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_21 = 0.064184
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21 = 0.17138
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_21 = -0.0010658
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21 = 0.02257
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_21 = 3.6971e-5
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_21 = 1.0823e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 022, W = 5.0u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_22 = 1.2591e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_22 = 7.8826e-20
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_22 = 0.016777
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22 = -26705.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22 = -0.13788
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_22 = 0.00085841
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22 = 0.032732
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_22 = -0.014452
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 023, W = 5.0u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_23 = -0.010788
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_23 = 3.3564e-11
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_23 = 3.011e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_23 = 0.00046251
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23 = 2290.4
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23 = 0.09276
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_23 = 0.00089335
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23 = 0.02941
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 024, W = 5.0u, L = 0.25u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24 = 0.084105
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_24 = 0.00034703
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24 = -0.027367
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_24 = -0.0082625
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_24 = 1.545e-11
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_24 = 2.4497e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_24 = -0.019165
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24 = -2665.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 025, W = 5.0u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25 = 34633.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25 = -0.49988
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_25 = 0.0009351
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25 = -0.014583
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_25 = -0.01222
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_25 = -1.5818e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_25 = 5.2715e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_25 = -0.01793
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_25 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 026, W = 7.0u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26 = 0.065303
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_26 = 0.00052886
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26 = -0.013059
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_26 = -0.0088359
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_26 = -5.3351e-11
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_26 = 1.8475e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_26 = -0.026142
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_26 = 0.022113
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_26 = -0.029735
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_26 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 027, W = 7.0u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27 = -0.044622
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_27 = -0.0004791
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27 = 0.014685
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_27 = 0.00017502
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_27 = 7.9422e-11
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_27 = -2.018e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_27 = 0.0050269
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_27 = -0.062963
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_27 = 0.073551
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 028, W = 7.0u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28 = 0.29531
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_28 = -0.0013902
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28 = 0.026712
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_28 = 0.0021134
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_28 = 1.9527e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_28 = -5.0295e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_28 = 0.020482
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_28 = -0.12263
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_28 = 0.068237
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 029, W = 7.0u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_29 = -0.11748
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_29 = 0.097986
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29 = 0.32486
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_29 = -0.0010323
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29 = 0.023278
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_29 = 2.5278e-5
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_29 = 1.7065e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_29 = -4.0984e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_29 = 0.019772
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 030, W = 7.0u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_30 = 0.0045478
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30 = -21113.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30 = 0.42541
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_30 = 0.0019309
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30 = 0.024852
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_30 = -0.030002
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_30 = 3.916e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_30 = -5.5528e-20
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 031, W = 7.0u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_31 = -0.026048
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31 = 11802.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31 = 0.057075
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_31 = 0.00062518
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31 = 0.00020745
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_31 = -0.016511
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_31 = -8.2694e-11
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_31 = 3.8486e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 032, W = 7.0u, L = 0.25u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_32 = 1.4441e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_32 = -0.021942
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32 = -3470.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32 = 0.10206
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_32 = 4.1162e-5
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32 = -0.020217
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_32 = -0.0072879
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_32 = 2.3274e-11
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 033, W = 7.0u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_33 = 4.3313e-12
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_33 = -3.3895e-20
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_33 = -0.0013118
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33 = 20.656
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33 = 0.60582
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_33 = -6.7689e-5
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33 = -0.015116
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_33 = 1.0469e-33
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 034, W = 0.42u, L = 1.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_34 = 0.022876
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_34 = 2.3669e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_34 = -2.6496e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_34 = 0.013143
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_34 = -1.7673e-8
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_34 = -5.2005e-9
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34 = -0.27625
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_34 = -0.0002157
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34 = -0.0097079
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 035, W = 0.42u, L = 20.0u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35 = 0.068952
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_35 = 0.00040549
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35 = -0.049997
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_35 = 0.0049572
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_35 = -1.1638e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_35 = 1.7782e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_35 = -0.0082316
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_35 = 2.7422e-8
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_35 = -3.9995e-9
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 036, W = 0.42u, L = 2.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36 = -39.498
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36 = 0.046265
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_36 = 0.00088129
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36 = -0.060841
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_36 = 0.0059014
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_36 = 2.124e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_36 = -1.0049e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_36 = -0.021848
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_36 = -7.7669e-8
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_36 = 2.8952e-8
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 037, W = 0.42u, L = 4.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_37 = -2.4687e-9
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37 = 0.0575
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_37 = 0.0036928
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37 = -0.078423
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_37 = -0.0036523
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_37 = -3.3052e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_37 = 1.3732e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_37 = -0.044816
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_37 = -1.2216e-7
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_37 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 038, W = 0.42u, L = 8.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_38 = -7.6337e-8
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_38 = 3.0215e-10
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38 = 0.056948
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_38 = 0.000428
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38 = -0.065945
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_38 = -0.0060343
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_38 = -5.9148e-11
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_38 = 1.5095e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_38 = -0.039769
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 039, W = 0.42u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39 = -0.016965
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_39 = -0.00027103
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39 = -7377.5
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39 = 0.022729
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_39 = -0.0032761
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_39 = 2.1113e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_39 = -3.3743e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_39 = 0.0068733
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_39 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 040, W = 0.42u, L = 0.18u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40 = 16736.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40 = -0.087082
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_40 = -0.0016136
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40 = 0.02991
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_40 = 0.00051508
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_40 = -5.6434e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_40 = 4.4059e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_40 = 0.038681
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_40 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 041, W = 0.42u, L = 0.5u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_41 = 0.036001
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41 = -18950.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41 = -0.1458
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_41 = -0.0010505
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41 = 0.032157
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_41 = 0.019753
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_41 = 1.3095e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_41 = -3.4743e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 042, W = 0.55u, L = 1.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_42 = -0.055461
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_42 = -1.9112e-7
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_42 = 9.0698e-11
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42 = 0.25017
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_42 = 0.0029063
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42 = -0.074951
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_42 = -0.011704
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_42 = -8.7192e-11
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_42 = 9.152e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 043, W = 0.55u, L = 2.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_43 = 1.0804e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_43 = -0.038517
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_43 = -1.0106e-7
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_43 = -3.2887e-9
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43 = 0.24291
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_43 = 0.0024377
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43 = -0.050427
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_43 = -0.0033063
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_43 = -1.8802e-10
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 044, W = 0.55u, L = 4.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_44 = -2.4438e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_44 = 1.0742e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_44 = -0.04155
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_44 = -1.4796e-7
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_44 = -3.1696e-9
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44 = 0.25082
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_44 = 0.0027361
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44 = -0.054247
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_44 = -0.0043806
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 045, W = 0.55u, L = 8.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_45 = -0.0079756
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_45 = -3.0833e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_45 = 1.0427e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_45 = -0.040223
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_45 = -1.1819e-7
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_45 = 1.8309e-10
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45 = 0.17754
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_45 = 0.0024422
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45 = -0.053285
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 046, W = 0.55u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46 = -0.22504
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_46 = -0.00091692
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46 = 0.0062628
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_46 = -0.015028
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_46 = -3.4e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_46 = 3.0008e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_46 = 0.043465
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46 = 70059.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 047, W = 0.55u, L = 0.5u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47 = -6190.8
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47 = -0.41079
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_47 = -0.00092357
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47 = -0.010036
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_47 = 0.0035187
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_47 = 3.1208e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_47 = -5.6959e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_47 = 0.0058894
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_47 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 048, W = 0.64u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48 = -7598.6
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48 = 0.059878
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_48 = -0.00011448
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48 = 0.014085
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_48 = -0.0060388
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_48 = 9.0006e-11
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_48 = -1.5016e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_48 = -0.0096942
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_48 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 049, W = 0.84u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49 = -10223.0
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49 = 0.21475
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_49 = 0.0030696
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49 = 0.041291
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_49 = -0.019245
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_49 = 1.4207e-9
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_49 = -1.3252e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_49 = -0.026095
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 050, W = 0.64u, L = 0.18u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50 = -13020.19512796
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_50 = -8.25379e-5
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50 = -0.74619177
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50 = -0.003959
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_50 = 0.00237687
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_50 = 1.76727e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_50 = -3.0963e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_50 = 0.08256679
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 051, W = 2.0u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51 = -13801.03896135
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_51 = 0.00045065
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51 = -0.33252405
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51 = 0.01885897
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_51 = 0.00023295
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_51 = 8.6482e-11
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_51 = 4.4521e-20
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_51 = 0.0486194
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_51 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 052, W = 1.12u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_52 = 0.05361098
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_52 = 1.83449e-7
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52 = -2407.39392921
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_52 = -0.00024377
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52 = -0.5622001
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52 = 0.00718778
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_52 = -0.001625
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_52 = -5.08997e-12
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_52 = -5.52904e-21
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 053, W = 1.65u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_53 = 0.06061
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53 = -21921.18384543
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_53 = 0.0002587
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53 = -0.32147005
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53 = 0.02092406
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_53 = 0.00113997
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_53 = 7.002e-11
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_53 = 1.26996e-21
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 054, W = 0.84u, L = 0.18u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_54 = -1.40124e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_54 = 0.02290802
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54 = -4076.48882566
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_54 = 0.00287678
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54 = -1.19974971
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54 = -0.00687001
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_54 = -0.009055
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_54 = 1.42864e-9
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 055, W = 1.68u, L = 0.18u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_55 = 1.94065e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_55 = -5.907e-20
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_55 = 0.03055499
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55 = -22283.99670468
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_55 = 0.00072546
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55 = 0.23037004
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55 = 0.01624287
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_55 = -0.00600001
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 056, W = 0.36u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_56 = -0.026
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56 = -7744.3
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_56 = -2.1326e-5
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56 = -0.040606
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 057, W = 0.54u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_57 = -0.00039634
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57 = -0.023293
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_57 = -0.021038
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_57 = -8.112e-8
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_57 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57 = 152000.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 058, W = 0.63u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58 = 78825.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_58 = -0.00031572
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58 = -0.0088034
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_58 = -0.021882
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_58 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_58 = -3.6053e-8
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_58 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 059, W = 0.7u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_59 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59 = 100000.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59 = -0.00118062
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_59 = 0.00058467
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59 = -0.90770424
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59 = -0.004599
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_59 = -0.021992
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_59 = 6.35098e-10
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_59 = -7.09206e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59 = 0.00022005
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_59 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_59 = 0.001118
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_59 = 0.06092346
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59 = -3.51778e-12
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_59 = 5.81762e-5
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_59 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 060, W = 0.75u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_60 = 5.92226e-5
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60 = 100000.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_60 = 0.0013154
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60 = -0.00120185
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60 = -1.02378836
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60 = -0.0049437
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_60 = -0.023394
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_60 = 9.55739e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_60 = -9.88789e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60 = 0.000224
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_60 = 0.04564715
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_60 = 0.0011381
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60 = -3.58105e-12
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 061, W = 0.79u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61 = -2.43054e-12
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_61 = 4.01958e-5
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_61 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_61 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61 = 484410.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61 = -0.00081573
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_61 = 0.0016786
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61 = -1.10667404
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61 = -0.0052213
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_61 = -0.02357
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_61 = 1.18041e-9
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_61 = -1.18473e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61 = 0.00015204
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_61 = 0.03487521
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_61 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_61 = 0.00077246
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 062, W = 0.82u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62 = -1.07843e-12
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_62 = 1.78349e-5
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62 = 442400.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62 = -0.00036194
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_62 = 0.0020028
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62 = -1.16381151
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62 = -0.0013335
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_62 = -0.022866
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_62 = 1.33329e-9
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_62 = -1.31807e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62 = 6.74589e-5
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_62 = 0.02751291
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_62 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_62 = 0.00034274
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 063, W = 0.82u, L = 0.18u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_63 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_63 = 0.00034274
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_63 = 0.02751293
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63 = -1.07843e-12
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_63 = 1.7835e-5
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_63 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_63 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63 = 100000.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63 = -0.00036194
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_63 = 0.0021034
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63 = -1.16381122
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63 = -0.00025003
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_63 = -0.014058
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_63 = 1.33329e-9
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_63 = -1.31807e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63 = 6.7459e-5
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 064, W = 0.82u, L = 0.25u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64 = 9.26987e-5
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64 = 348355.7500906
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_64 = 0.00037141
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_64 = -0.00038001
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_64 = 0.02171056
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64 = -1.25142e-12
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_64 = -2.77702e-5
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_64 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_64 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64 = 31804.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_64 = -0.00054783
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64 = -0.17599174
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64 = -0.025021
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_64 = -0.014998
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_64 = 4.72444e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_64 = -7.42909e-19
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 065, W = 0.82u, L = 0.5u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65 = 50000.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_65 = -0.00079087
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65 = -0.026825
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_65 = -0.0094836
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_65 = 0.0
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 066, W = 0.86u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_66 = 1.21828e-9
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_66 = -1.19646e-18
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_66 = -0.00025474
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_66 = 0.0273647
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66 = 3.61331e-13
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_66 = -1.52588e-6
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66 = 484680.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_66 = 0.0017686
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66 = -1.10730207
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66 = 0.0028658
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_66 = -0.022338
*
* sky130_fd_pr__pfet_01v8_hvt, Bin 067, W = 0.94u, L = 0.15u
* ------------------------------------
+ sky130_fd_pr__pfet_01v8_hvt__k2_diff_67 = -0.0168
+ sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ua_diff_67 = 4.71861e-10
+ sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ub_diff_67 = -4.69835e-19
+ sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67 = -6.2769e-5
+ sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__ags_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__a0_diff_67 = -0.00045296
+ sky130_fd_pr__pfet_01v8_hvt__voff_diff_67 = 0.04331183
+ sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67 = 6.42491e-13
+ sky130_fd_pr__pfet_01v8_hvt__keta_diff_67 = -2.71304e-6
+ sky130_fd_pr__pfet_01v8_hvt__b0_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__b1_diff_67 = 0.0
+ sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67 = 500000.0
+ sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67 = -3.68096e-5
+ sky130_fd_pr__pfet_01v8_hvt__u0_diff_67 = 0.00028484
+ sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67 = -0.77623339
+ sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67 = 0.012571
*.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8_hvt.pm3.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8_hvt__ss.pm3.spice"
