* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 38
.param
+ sky130_fd_pr__nfet_01v8_lvt__toxe_mult = 0.9635
+ sky130_fd_pr__nfet_01v8_lvt__rshn_mult = 1.0
+ sky130_fd_pr__nfet_01v8_lvt__overlap_mult = 0.88119
+ sky130_fd_pr__nfet_01v8_lvt__ajunction_mult = 0.87784
+ sky130_fd_pr__nfet_01v8_lvt__pjunction_mult = 0.78244
+ sky130_fd_pr__nfet_01v8_lvt__lint_diff = 1.21275e-8
+ sky130_fd_pr__nfet_01v8_lvt__wint_diff = -2.252e-8
+ sky130_fd_pr__nfet_01v8_lvt__dlc_diff = 7.7131e-9
+ sky130_fd_pr__nfet_01v8_lvt__dwc_diff = -2.252e-8
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 000, W = 1.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_0 = -0.064001
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_0 = 0.0081134
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_0 = 0.0020103
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_0 = -0.10975
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_0 = -7.0587e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_0 = 3.8853e-19
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0 = 0.70456
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0 = -0.0076786
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 001, W = 1.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_1 = -0.050662
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_1 = 0.0077884
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_1 = -0.10908
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_1 = 0.00093901
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_1 = 6.8072e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_1 = 2.826e-19
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1 = 0.39852
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1 = -0.0078928
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 002, W = 1.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2 = -0.0043298
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_2 = 0.0090734
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_2 = 0.0099409
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_2 = -0.0061366
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_2 = 0.00062214
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_2 = -1.9272e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_2 = 2.575e-19
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2 = 0.72829
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 003, W = 1.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3 = 1.4729
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3 = -0.058087
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_3 = 0.031103
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_3 = -0.0015859
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_3 = 6.8273e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3 = -26072.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_3 = 1.612e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 004, W = 1.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4 = 1.5178
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4 = -0.082199
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_4 = 0.019857
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_4 = -0.0021861
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_4 = 1.8015e-11
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4 = -21912.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_4 = 4.5553e-20
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 005, W = 1.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_5 = 4.5063e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5 = 0.95603
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5 = -0.011184
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_5 = 0.0093294
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_5 = 0.0024348
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_5 = -2.0398e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5 = -12947.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_5 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 006, W = 1.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_6 = 2.7444e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6 = 1.3429
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6 = -0.010655
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_6 = -0.00062272
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_6 = 0.0005695
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_6 = -3.92e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6 = -10142.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_6 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 007, W = 3.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_7 = 2.4261e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7 = 0.77503
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7 = 8.7015e-5
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_7 = -0.026006
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_7 = 0.0038481
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_7 = -0.035935
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_7 = 0.0013497
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_7 = -2.3833e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 008, W = 3.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_8 = -0.034253
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_8 = 0.00070921
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_8 = -5.0806e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_8 = 1.9943e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8 = 0.36129
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8 = -0.0057838
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_8 = -0.020934
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_8 = 0.0013629
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 009, W = 3.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_9 = -0.006192
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_9 = 0.00026333
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_9 = -1.1842e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_9 = 1.3971e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9 = 0.42662
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9 = -0.00025391
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_9 = 0.0058881
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_9 = 0.0058275
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 010, W = 3.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_10 = 3.5409e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_10 = -1.1456e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_10 = -0.0028995
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10 = -19021.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10 = -0.085201
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10 = 1.2225
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_10 = 0.033776
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 011, W = 3.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_11 = 0.024793
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_11 = 2.1273e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_11 = 1.6509e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_11 = -0.00039822
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11 = -12938.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11 = -0.063158
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11 = 1.2006
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 012, W = 3.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_12 = 0.014212
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_12 = -8.5273e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_12 = 4.9607e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_12 = 0.0012429
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12 = -7928.4
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12 = -0.020197
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12 = 0.93234
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_12 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 013, W = 3.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_13 = 0.012015
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_13 = 9.2164e-14
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_13 = 2.3157e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_13 = 0.00020896
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13 = -6126.5
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13 = -0.0076636
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13 = 1.2266
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_13 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 014, W = 5.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14 = 0.63062
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_14 = 0.0029183
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_14 = -1.0862e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_14 = 2.207e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_14 = -0.033478
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_14 = -0.050039
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_14 = 0.00097848
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14 = -0.0082701
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 015, W = 5.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15 = 0.00092243
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15 = 0.51633
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_15 = -0.0060606
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_15 = -1.8742e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_15 = 2.3666e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_15 = 0.011196
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_15 = 0.015378
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_15 = 0.00093567
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 016, W = 5.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_16 = -0.02206
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_16 = 0.00051071
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16 = -0.010136
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16 = 0.10272
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_16 = 0.0085836
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_16 = 1.3225e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_16 = 1.6378e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_16 = 0.0031853
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 017, W = 5.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_17 = -0.00082717
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17 = -13818.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17 = -0.074175
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17 = 1.3395
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_17 = 0.037049
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_17 = 2.9203e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_17 = 1.1213e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 018, W = 5.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_18 = -0.0012159
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18 = -16297.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18 = -0.047066
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18 = 1.2712
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_18 = 0.025327
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_18 = 2.6552e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_18 = 8.029e-20
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 019, W = 5.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_19 = 3.6615e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_19 = 0.00042198
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19 = -13450.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19 = -0.028005
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19 = 0.75655
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_19 = 0.011293
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_19 = -3.8741e-11
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 020, W = 5.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_20 = -2.0719e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_20 = 2.5573e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_20 = 0.00081091
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20 = -899.91
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20 = -0.011093
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20 = 1.1478
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_20 = 0.0019437
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 021, W = 7.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_21 = -4.2056e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_21 = 2.5388e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_21 = 0.045409
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_21 = 0.048057
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_21 = 0.0013807
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21 = 0.00038533
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21 = 0.74534
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_21 = -0.0047384
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 022, W = 7.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_22 = 0.0076765
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_22 = -1.281e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_22 = 1.9584e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_22 = 0.00072066
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_22 = -0.0067956
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_22 = 0.00074354
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22 = -0.0053605
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22 = 0.45602
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 023, W = 7.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_23 = 0.0067583
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_23 = -2.3598e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_23 = 2.1315e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_23 = -0.00059699
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_23 = 0.031865
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_23 = 0.0010023
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23 = -0.004118
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23 = 0.3288
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_23 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 024, W = 7.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_24 = 0.038683
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_24 = 1.1967e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_24 = -1.6049e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_24 = -0.0047096
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24 = -14167.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24 = -0.089849
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24 = 1.3376
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_24 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 025, W = 7.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25 = 1.2419
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_25 = 0.022825
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_25 = 6.4936e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_25 = -2.5046e-21
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_25 = -0.0023153
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25 = -15924.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25 = -0.046521
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 026, W = 7.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26 = -0.018801
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26 = 0.73783
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_26 = 0.01227
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_26 = -1.2398e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_26 = 3.5666e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_26 = 0.0014372
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26 = -11322.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 027, W = 7.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_27 = 0.00066763
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27 = -1962.1
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27 = -0.0048024
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27 = 0.98774
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_27 = 0.0037101
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_27 = -2.8272e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_27 = 2.1671e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 028, W = 0.42u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_28 = 0.002882
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28 = -0.018416
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28 = 0.13245
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_28 = 9.6413e-8
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_28 = 1.0459e-9
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_28 = 0.0046606
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_28 = -1.7631e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_28 = 5.0687e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 029, W = 0.42u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_29 = -0.0019238
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29 = -26661.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29 = -0.11716
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29 = 1.6054
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_29 = 0.029703
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_29 = 4.346e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_29 = 1.5069e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 030, W = 0.42u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_30 = 6.8804e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_30 = -0.00058909
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30 = -22958.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30 = -0.10542
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30 = 1.5302
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_30 = 0.012433
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_30 = 2.2286e-11
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 031, W = 0.55u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_31 = 2.689e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_31 = -3.4876e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_31 = -0.0029007
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31 = -34751.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31 = -0.13397
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31 = 2.1416
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_31 = 0.017083
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 032, W = 0.64u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_32 = 2.0615e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_32 = 3.0798e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_32 = -0.0015571
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32 = -19624.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32 = -0.13512
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32 = 2.159
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_32 = 0.017306
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 033, W = 0.84u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_33 = 0.016181
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_33 = 2.0951e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_33 = -7.6709e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_33 = -0.0019419
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33 = -15572.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33 = -0.12569
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33 = 1.9124
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 034, W = 1.65u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_34 = 0.031783
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_34 = 1.2373e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_34 = -1.044e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_34 = -0.0033755
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34 = -17260.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34 = -0.087483
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34 = 1.646
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_34 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 035, W = 3.01u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_35 = 0.032894
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_35 = 2.3003e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_35 = -7.6801e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_35 = -0.0030264
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35 = -21178.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35 = -0.083109
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35 = 1.2691
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_35 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 036, W = 5.05u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36 = 1.4374
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_36 = 0.037302
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_36 = 9.319e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_36 = 1.7106e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_36 = -0.00099139
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36 = -13868.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36 = -0.071658
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 037, W = 5.05u, L = 0.25u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37 = -0.023221
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37 = 0.89187
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_37 = 0.010877
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_37 = -2.1819e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_37 = 3.2503e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_37 = 0.00072118
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37 = -12287.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_01v8_lvt.pm3.spice"
