* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 52
.param
+ sky130_fd_pr__pfet_01v8__toxe_mult = 0.9635
+ sky130_fd_pr__pfet_01v8__rshp_mult = 1.0
+ sky130_fd_pr__pfet_01v8__overlap_mult = 0.88516
+ sky130_fd_pr__pfet_01v8__ajunction_mult = 0.93001
+ sky130_fd_pr__pfet_01v8__pjunction_mult = 0.93439
+ sky130_fd_pr__pfet_01v8__lint_diff = 1.21275e-8
+ sky130_fd_pr__pfet_01v8__wint_diff = -2.252e-8
+ sky130_fd_pr__pfet_01v8__dlc_diff = 1.21275e-8
+ sky130_fd_pr__pfet_01v8__dwc_diff = -2.252e-8
*
* sky130_fd_pr__pfet_01v8, Bin 000, W = 1.26u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_0 = 1.986
+ sky130_fd_pr__pfet_01v8__vsat_diff_0 = 2943.9
+ sky130_fd_pr__pfet_01v8__a0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_0 = -8.9653e-12
+ sky130_fd_pr__pfet_01v8__keta_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_0 = -0.0060133
+ sky130_fd_pr__pfet_01v8__vth0_diff_0 = -0.015634
+ sky130_fd_pr__pfet_01v8__pditsd_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_0 = 0.00062824
+ sky130_fd_pr__pfet_01v8__b1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_0 = -0.20331
+ sky130_fd_pr__pfet_01v8__ags_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_0 = 3.0962e-19
*
* sky130_fd_pr__pfet_01v8, Bin 001, W = 1.68u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_1 = 2.3976e-19
+ sky130_fd_pr__pfet_01v8__agidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_1 = 1.9897
+ sky130_fd_pr__pfet_01v8__vsat_diff_1 = -5832.9
+ sky130_fd_pr__pfet_01v8__a0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_1 = -5.1977e-11
+ sky130_fd_pr__pfet_01v8__keta_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_1 = -0.0097727
+ sky130_fd_pr__pfet_01v8__vth0_diff_1 = -0.079534
+ sky130_fd_pr__pfet_01v8__pditsd_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_1 = 0.00032864
+ sky130_fd_pr__pfet_01v8__b1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_1 = -0.18643
+ sky130_fd_pr__pfet_01v8__ags_diff_1 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 002, W = 1.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_2 = -0.096547
+ sky130_fd_pr__pfet_01v8__ags_diff_2 = 0.14368
+ sky130_fd_pr__pfet_01v8__bgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_2 = 4.385e-19
+ sky130_fd_pr__pfet_01v8__agidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_2 = -0.19028
+ sky130_fd_pr__pfet_01v8__vsat_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_2 = -0.1314
+ sky130_fd_pr__pfet_01v8__pdits_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_2 = -2.3189e-11
+ sky130_fd_pr__pfet_01v8__keta_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_2 = -0.0084567
+ sky130_fd_pr__pfet_01v8__vth0_diff_2 = 0.0096478
+ sky130_fd_pr__pfet_01v8__pditsd_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_2 = 0.002096
+ sky130_fd_pr__pfet_01v8__b1_diff_2 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 003, W = 1.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__b1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_3 = -0.091929
+ sky130_fd_pr__pfet_01v8__ags_diff_3 = 0.044206
+ sky130_fd_pr__pfet_01v8__bgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_3 = 5.1919e-19
+ sky130_fd_pr__pfet_01v8__nfactor_diff_3 = 0.10772
+ sky130_fd_pr__pfet_01v8__vsat_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_3 = -0.048991
+ sky130_fd_pr__pfet_01v8__pdits_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_3 = -5.7469e-12
+ sky130_fd_pr__pfet_01v8__keta_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_3 = -0.012618
+ sky130_fd_pr__pfet_01v8__vth0_diff_3 = 0.01485
+ sky130_fd_pr__pfet_01v8__pditsd_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_3 = 0.0026341
*
* sky130_fd_pr__pfet_01v8, Bin 004, W = 1.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_4 = 0.0026249
+ sky130_fd_pr__pfet_01v8__vth0_diff_4 = 0.00098819
+ sky130_fd_pr__pfet_01v8__b1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_4 = -0.091492
+ sky130_fd_pr__pfet_01v8__ags_diff_4 = 0.044861
+ sky130_fd_pr__pfet_01v8__ub_diff_4 = 4.9172e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_4 = 0.10992
+ sky130_fd_pr__pfet_01v8__vsat_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_4 = -0.044825
+ sky130_fd_pr__pfet_01v8__pdits_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_4 = -3.8288e-12
+ sky130_fd_pr__pfet_01v8__keta_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_4 = -0.013534
*
* sky130_fd_pr__pfet_01v8, Bin 005, W = 1.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__keta_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_5 = -0.01509
+ sky130_fd_pr__pfet_01v8__pditsd_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_5 = 0.0021952
+ sky130_fd_pr__pfet_01v8__vth0_diff_5 = -0.013252
+ sky130_fd_pr__pfet_01v8__b1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_5 = -0.10553
+ sky130_fd_pr__pfet_01v8__cgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_5 = 0.082407
+ sky130_fd_pr__pfet_01v8__ub_diff_5 = 4.3295e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_5 = 0.16171
+ sky130_fd_pr__pfet_01v8__vsat_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_5 = -0.077052
+ sky130_fd_pr__pfet_01v8__pdits_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_5 = -1.4191e-11
+ sky130_fd_pr__pfet_01v8__rdsw_diff_5 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 006, W = 1.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_6 = -1.0000e-2
+ sky130_fd_pr__pfet_01v8__pditsd_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_6 = -2.9577e-4
+ sky130_fd_pr__pfet_01v8__vth0_diff_6 = -9.0696e-2
+ sky130_fd_pr__pfet_01v8__b1_diff_6 = 8.2483e-11
+ sky130_fd_pr__pfet_01v8__voff_diff_6 = -0.17179
+ sky130_fd_pr__pfet_01v8__cgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_6 = 7.825e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_6 = 1.8740
+ sky130_fd_pr__pfet_01v8__vsat_diff_6 = -10439.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_6 = -4.9969e-10
+ sky130_fd_pr__pfet_01v8__pclm_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_6 = -4.8816e-10
*
* sky130_fd_pr__pfet_01v8, Bin 007, W = 1.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_7 = -2.0991e-12
+ sky130_fd_pr__pfet_01v8__rdsw_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_7 = -0.0065174
+ sky130_fd_pr__pfet_01v8__pditsd_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_7 = 0.00043857
+ sky130_fd_pr__pfet_01v8__vth0_diff_7 = -0.062759
+ sky130_fd_pr__pfet_01v8__b1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_7 = -0.24284
+ sky130_fd_pr__pfet_01v8__cgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_7 = 2.367e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_7 = 1.4003
+ sky130_fd_pr__pfet_01v8__vsat_diff_7 = -5947.7
+ sky130_fd_pr__pfet_01v8__agidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_7 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 008, W = 1.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_8 = 3.035e-12
+ sky130_fd_pr__pfet_01v8__rdsw_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_8 = -0.004591
+ sky130_fd_pr__pfet_01v8__pditsd_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_8 = 1.433e-5
+ sky130_fd_pr__pfet_01v8__vth0_diff_8 = 0.028589
+ sky130_fd_pr__pfet_01v8__b1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_8 = -0.1765
+ sky130_fd_pr__pfet_01v8__cgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_8 = 2.1102e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_8 = 0.61687
+ sky130_fd_pr__pfet_01v8__vsat_diff_8 = 24692.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_8 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 009, W = 1.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_9 = -4.8794e-12
+ sky130_fd_pr__pfet_01v8__rdsw_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_9 = -0.0092108
+ sky130_fd_pr__pfet_01v8__pditsd_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_9 = 0.0011423
+ sky130_fd_pr__pfet_01v8__vth0_diff_9 = 0.038262
+ sky130_fd_pr__pfet_01v8__b1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_9 = -0.097594
+ sky130_fd_pr__pfet_01v8__cgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_9 = 3.4941e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_9 = 0.089772
+ sky130_fd_pr__pfet_01v8__vsat_diff_9 = 15016.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_9 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 010, W = 2.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_10 = -12128.0
+ sky130_fd_pr__pfet_01v8__u0_diff_10 = -0.00052194
+ sky130_fd_pr__pfet_01v8__vth0_diff_10 = -0.052713
+ sky130_fd_pr__pfet_01v8__cgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_10 = -2.3474e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_10 = 0.79321
+ sky130_fd_pr__pfet_01v8__ub_diff_10 = 2.4004e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_10 = 0.024155
+ sky130_fd_pr__pfet_01v8__voff_diff_10 = -0.12071
+ sky130_fd_pr__pfet_01v8__a0_diff_10 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 011, W = 3.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_11 = -0.090266
+ sky130_fd_pr__pfet_01v8__a0_diff_11 = -0.13175
+ sky130_fd_pr__pfet_01v8__pditsd_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_11 = 31999.0
+ sky130_fd_pr__pfet_01v8__u0_diff_11 = 0.001628
+ sky130_fd_pr__pfet_01v8__vth0_diff_11 = -0.00098349
+ sky130_fd_pr__pfet_01v8__cgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_11 = -4.1402e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_11 = 0.078308
+ sky130_fd_pr__pfet_01v8__ub_diff_11 = 4.0944e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_11 = 0.10901
+ sky130_fd_pr__pfet_01v8__k2_diff_11 = -0.014602
*
* sky130_fd_pr__pfet_01v8, Bin 012, W = 3.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_12 = 0.10005
+ sky130_fd_pr__pfet_01v8__k2_diff_12 = -0.0086498
+ sky130_fd_pr__pfet_01v8__voff_diff_12 = -0.085532
+ sky130_fd_pr__pfet_01v8__a0_diff_12 = -0.11393
+ sky130_fd_pr__pfet_01v8__pditsd_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_12 = 0.0020542
+ sky130_fd_pr__pfet_01v8__vth0_diff_12 = 0.00065633
+ sky130_fd_pr__pfet_01v8__cgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_12 = -9.5084e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_12 = 0.057478
+ sky130_fd_pr__pfet_01v8__ub_diff_12 = 4.1587e-19
*
* sky130_fd_pr__pfet_01v8, Bin 013, W = 3.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_13 = 0.095358
+ sky130_fd_pr__pfet_01v8__ub_diff_13 = 4.1151e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_13 = 0.05372
+ sky130_fd_pr__pfet_01v8__k2_diff_13 = -0.00679
+ sky130_fd_pr__pfet_01v8__voff_diff_13 = -0.075626
+ sky130_fd_pr__pfet_01v8__a0_diff_13 = -0.060887
+ sky130_fd_pr__pfet_01v8__eta0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_13 = 0.0021092
+ sky130_fd_pr__pfet_01v8__vsat_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_13 = 0.010222
+ sky130_fd_pr__pfet_01v8__cgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_13 = -3.3811e-12
*
* sky130_fd_pr__pfet_01v8, Bin 014, W = 3.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_14 = -1.9824e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_14 = 0.025266
+ sky130_fd_pr__pfet_01v8__ub_diff_14 = 4.9458e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_14 = 0.012252
+ sky130_fd_pr__pfet_01v8__k2_diff_14 = -0.0067467
+ sky130_fd_pr__pfet_01v8__voff_diff_14 = -0.072864
+ sky130_fd_pr__pfet_01v8__eta0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_14 = -0.067604
+ sky130_fd_pr__pfet_01v8__pditsd_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_14 = 0.002432
+ sky130_fd_pr__pfet_01v8__vsat_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_14 = 0.012639
+ sky130_fd_pr__pfet_01v8__cgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_14 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 015, W = 3.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_15 = -3.1715e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_15 = 1.8982
+ sky130_fd_pr__pfet_01v8__ub_diff_15 = 1.5817e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_15 = -0.0056566
+ sky130_fd_pr__pfet_01v8__pdits_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_15 = -0.152
+ sky130_fd_pr__pfet_01v8__eta0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_15 = 0.00027437
+ sky130_fd_pr__pfet_01v8__vsat_diff_15 = -11954.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_15 = -0.10163
+ sky130_fd_pr__pfet_01v8__cgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_15 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 016, W = 3.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_16 = 2.484e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_16 = 1.065
+ sky130_fd_pr__pfet_01v8__tvoff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_16 = 1.6562e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_16 = -0.004036
+ sky130_fd_pr__pfet_01v8__pdits_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_16 = -0.23592
+ sky130_fd_pr__pfet_01v8__eta0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_16 = 0.00046849
+ sky130_fd_pr__pfet_01v8__vsat_diff_16 = -1875.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_16 = -0.048685
+ sky130_fd_pr__pfet_01v8__cgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_16 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 017, W = 3.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_17 = 0.4592
+ sky130_fd_pr__pfet_01v8__ua_diff_17 = -4.9962e-11
+ sky130_fd_pr__pfet_01v8__tvoff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_17 = 2.2716e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_17 = -0.00074906
+ sky130_fd_pr__pfet_01v8__pdits_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_17 = -0.17242
+ sky130_fd_pr__pfet_01v8__eta0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_17 = 0.00022565
+ sky130_fd_pr__pfet_01v8__vsat_diff_17 = 60423.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_17 = -0.024518
+ sky130_fd_pr__pfet_01v8__cgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_17 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 018, W = 3.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_18 = 0.31736
+ sky130_fd_pr__pfet_01v8__ua_diff_18 = -3.6007e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_18 = 2.7771e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_18 = -0.013233
+ sky130_fd_pr__pfet_01v8__pdits_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_18 = -0.11303
+ sky130_fd_pr__pfet_01v8__eta0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_18 = 0.0012188
+ sky130_fd_pr__pfet_01v8__vsat_diff_18 = 43395.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_18 = 0.014578
+ sky130_fd_pr__pfet_01v8__cgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_18 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 019, W = 5.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_19 = -0.25759
+ sky130_fd_pr__pfet_01v8__ua_diff_19 = -3.3858e-11
+ sky130_fd_pr__pfet_01v8__tvoff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_19 = 0.18403
+ sky130_fd_pr__pfet_01v8__ub_diff_19 = 2.7193e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_19 = -0.0095727
+ sky130_fd_pr__pfet_01v8__pdits_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_19 = -0.08029
+ sky130_fd_pr__pfet_01v8__eta0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_19 = -0.18799
+ sky130_fd_pr__pfet_01v8__pditsd_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_19 = 0.0011002
+ sky130_fd_pr__pfet_01v8__vsat_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_19 = 0.01782
*
* sky130_fd_pr__pfet_01v8, Bin 020, W = 5.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__u0_diff_20 = 0.0013275
+ sky130_fd_pr__pfet_01v8__vth0_diff_20 = 0.013401
+ sky130_fd_pr__pfet_01v8__cgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_20 = -3.6861e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_20 = 0.10548
+ sky130_fd_pr__pfet_01v8__ub_diff_20 = 2.5181e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_20 = 0.048702
+ sky130_fd_pr__pfet_01v8__k2_diff_20 = -0.0096983
+ sky130_fd_pr__pfet_01v8__voff_diff_20 = -0.069333
+ sky130_fd_pr__pfet_01v8__a0_diff_20 = -0.054389
+ sky130_fd_pr__pfet_01v8__pditsd_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_20 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 021, W = 5.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_21 = 0.0017616
+ sky130_fd_pr__pfet_01v8__vth0_diff_21 = 0.016691
+ sky130_fd_pr__pfet_01v8__cgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_21 = -3.2379e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_21 = 0.097273
+ sky130_fd_pr__pfet_01v8__ub_diff_21 = 3.1768e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_21 = 0.039634
+ sky130_fd_pr__pfet_01v8__k2_diff_21 = -0.010143
+ sky130_fd_pr__pfet_01v8__voff_diff_21 = -0.065522
+ sky130_fd_pr__pfet_01v8__a0_diff_21 = -0.042736
*
* sky130_fd_pr__pfet_01v8, Bin 022, W = 5.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_22 = -0.065062
+ sky130_fd_pr__pfet_01v8__a0_diff_22 = -0.04183
+ sky130_fd_pr__pfet_01v8__pditsd_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_22 = 0.0019576
+ sky130_fd_pr__pfet_01v8__vth0_diff_22 = 0.011363
+ sky130_fd_pr__pfet_01v8__cgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_22 = -3.3906e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_22 = 0.1184
+ sky130_fd_pr__pfet_01v8__ub_diff_22 = 3.5796e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_22 = 0.037149
+ sky130_fd_pr__pfet_01v8__k2_diff_22 = -0.010219
*
* sky130_fd_pr__pfet_01v8, Bin 023, W = 5.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_23 = -0.0010754
+ sky130_fd_pr__pfet_01v8__voff_diff_23 = -0.18456
+ sky130_fd_pr__pfet_01v8__a0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_23 = -8584.1
+ sky130_fd_pr__pfet_01v8__u0_diff_23 = 9.6021e-5
+ sky130_fd_pr__pfet_01v8__vth0_diff_23 = -0.10786
+ sky130_fd_pr__pfet_01v8__cgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_23 = -6.7208e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_23 = 1.5227
+ sky130_fd_pr__pfet_01v8__ub_diff_23 = 1.6075e-19
*
* sky130_fd_pr__pfet_01v8, Bin 024, W = 5.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_24 = 1.0638
+ sky130_fd_pr__pfet_01v8__ub_diff_24 = 1.1879e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_24 = -0.00089499
+ sky130_fd_pr__pfet_01v8__voff_diff_24 = -0.212
+ sky130_fd_pr__pfet_01v8__a0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_24 = 0.00015187
+ sky130_fd_pr__pfet_01v8__vsat_diff_24 = 10165.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_24 = -0.060941
+ sky130_fd_pr__pfet_01v8__cgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_24 = -1.8608e-11
*
* sky130_fd_pr__pfet_01v8, Bin 025, W = 5.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_25 = -7.047e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_25 = 0.31553
+ sky130_fd_pr__pfet_01v8__ub_diff_25 = 1.7579e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_25 = -0.002567
+ sky130_fd_pr__pfet_01v8__voff_diff_25 = -0.14026
+ sky130_fd_pr__pfet_01v8__eta0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_25 = 0.00048574
+ sky130_fd_pr__pfet_01v8__vsat_diff_25 = 17176.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_25 = -0.03724
+ sky130_fd_pr__pfet_01v8__cgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_25 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 026, W = 5.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_26 = 8.7232e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_26 = 0.26077
+ sky130_fd_pr__pfet_01v8__ub_diff_26 = 2.6738e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_26 = -0.012506
+ sky130_fd_pr__pfet_01v8__pdits_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_26 = -0.078182
+ sky130_fd_pr__pfet_01v8__eta0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_26 = 0.0013823
+ sky130_fd_pr__pfet_01v8__vsat_diff_26 = 5999.4
+ sky130_fd_pr__pfet_01v8__vth0_diff_26 = 0.0080947
+ sky130_fd_pr__pfet_01v8__cgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_26 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 027, W = 7.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_27 = -1.4834e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_27 = -0.083423
+ sky130_fd_pr__pfet_01v8__tvoff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_27 = 0.1249
+ sky130_fd_pr__pfet_01v8__ub_diff_27 = 2.9424e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_27 = -0.0086855
+ sky130_fd_pr__pfet_01v8__pdits_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_27 = -0.059765
+ sky130_fd_pr__pfet_01v8__eta0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_27 = -0.1799
+ sky130_fd_pr__pfet_01v8__pditsd_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_27 = 0.0013548
+ sky130_fd_pr__pfet_01v8__vsat_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_27 = 0.0081694
+ sky130_fd_pr__pfet_01v8__cgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_27 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 028, W = 7.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_28 = 0.033842
+ sky130_fd_pr__pfet_01v8__ua_diff_28 = -9.0908e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_28 = 0.093633
+ sky130_fd_pr__pfet_01v8__ub_diff_28 = 2.7565e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_28 = -0.011195
+ sky130_fd_pr__pfet_01v8__pdits_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_28 = -0.065187
+ sky130_fd_pr__pfet_01v8__eta0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_28 = -0.10433
+ sky130_fd_pr__pfet_01v8__pditsd_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_28 = 0.0014348
+ sky130_fd_pr__pfet_01v8__vsat_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_28 = 0.015055
+ sky130_fd_pr__pfet_01v8__cgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_28 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 029, W = 7.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_29 = 0.10459
+ sky130_fd_pr__pfet_01v8__ua_diff_29 = -3.8377e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_29 = 0.044466
+ sky130_fd_pr__pfet_01v8__ub_diff_29 = 3.6296e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_29 = -0.010687
+ sky130_fd_pr__pfet_01v8__pdits_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_29 = -0.067361
+ sky130_fd_pr__pfet_01v8__eta0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_29 = -0.052347
+ sky130_fd_pr__pfet_01v8__pditsd_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_29 = 0.0020174
+ sky130_fd_pr__pfet_01v8__vsat_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_29 = 0.011199
+ sky130_fd_pr__pfet_01v8__cgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_29 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 030, W = 7.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_30 = -3.165e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_30 = 0.15193
+ sky130_fd_pr__pfet_01v8__ub_diff_30 = 3.9189e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_30 = 0.044301
+ sky130_fd_pr__pfet_01v8__k2_diff_30 = -0.011203
+ sky130_fd_pr__pfet_01v8__voff_diff_30 = -0.077571
+ sky130_fd_pr__pfet_01v8__a0_diff_30 = -0.048631
+ sky130_fd_pr__pfet_01v8__pditsd_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_30 = 0.0019907
+ sky130_fd_pr__pfet_01v8__vth0_diff_30 = 0.0094697
*
* sky130_fd_pr__pfet_01v8, Bin 031, W = 7.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__u0_diff_31 = 0.00011508
+ sky130_fd_pr__pfet_01v8__vth0_diff_31 = -0.10527
+ sky130_fd_pr__pfet_01v8__cgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_31 = -2.3155e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_31 = 1.2874
+ sky130_fd_pr__pfet_01v8__ub_diff_31 = 8.4151e-20
+ sky130_fd_pr__pfet_01v8__pdits_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_31 = -0.0058092
+ sky130_fd_pr__pfet_01v8__voff_diff_31 = -0.16551
+ sky130_fd_pr__pfet_01v8__a0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_31 = -7742.4
*
* sky130_fd_pr__pfet_01v8, Bin 032, W = 7.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_32 = 3510.8
+ sky130_fd_pr__pfet_01v8__u0_diff_32 = 0.00026428
+ sky130_fd_pr__pfet_01v8__vth0_diff_32 = -0.061382
+ sky130_fd_pr__pfet_01v8__cgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_32 = 1.8292e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_32 = 0.65166
+ sky130_fd_pr__pfet_01v8__ub_diff_32 = 9.7474e-20
+ sky130_fd_pr__pfet_01v8__pdits_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_32 = -0.0047382
+ sky130_fd_pr__pfet_01v8__voff_diff_32 = -0.12042
+ sky130_fd_pr__pfet_01v8__a0_diff_32 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 033, W = 7.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_33 = -0.096282
+ sky130_fd_pr__pfet_01v8__a0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_33 = 23751.0
+ sky130_fd_pr__pfet_01v8__u0_diff_33 = 0.00039004
+ sky130_fd_pr__pfet_01v8__vth0_diff_33 = -0.034284
+ sky130_fd_pr__pfet_01v8__cgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_33 = -1.7562e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_33 = 0.15621
+ sky130_fd_pr__pfet_01v8__ub_diff_33 = 1.6062e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_33 = -0.0052902
*
* sky130_fd_pr__pfet_01v8, Bin 034, W = 7.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_34 = -0.012412
+ sky130_fd_pr__pfet_01v8__voff_diff_34 = -0.07986
+ sky130_fd_pr__pfet_01v8__a0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_34 = 3998.9
+ sky130_fd_pr__pfet_01v8__u0_diff_34 = 0.0014177
+ sky130_fd_pr__pfet_01v8__vth0_diff_34 = 0.0026179
+ sky130_fd_pr__pfet_01v8__cgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_34 = 1.2144e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_34 = 0.2897
+ sky130_fd_pr__pfet_01v8__ub_diff_34 = 2.9051e-19
*
* sky130_fd_pr__pfet_01v8, Bin 035, W = 0.42u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_35 = 0.65595
+ sky130_fd_pr__pfet_01v8__ub_diff_35 = 4.9108e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_35 = -0.0082856
+ sky130_fd_pr__pfet_01v8__voff_diff_35 = -0.14486
+ sky130_fd_pr__pfet_01v8__a0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_35 = 0.0027403
+ sky130_fd_pr__pfet_01v8__vsat_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_35 = 0.00018011
+ sky130_fd_pr__pfet_01v8__cgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_35 = -2.68e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_35 = -3.7723e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_35 = 5.0827e-12
*
* sky130_fd_pr__pfet_01v8, Bin 036, W = 0.42u, L = 20.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_36 = 4.3216e-10
+ sky130_fd_pr__pfet_01v8__ua_diff_36 = -4.8976e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_36 = 0.29381
+ sky130_fd_pr__pfet_01v8__ub_diff_36 = 4.2986e-20
+ sky130_fd_pr__pfet_01v8__pdits_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_36 = -0.0015247
+ sky130_fd_pr__pfet_01v8__voff_diff_36 = -0.098227
+ sky130_fd_pr__pfet_01v8__eta0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_36 = 0.00017694
+ sky130_fd_pr__pfet_01v8__vsat_diff_36 = 20007.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_36 = 0.026332
+ sky130_fd_pr__pfet_01v8__cgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_36 = -5.3679e-8
*
* sky130_fd_pr__pfet_01v8, Bin 037, W = 0.42u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_37 = -5.8281e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_37 = 4.8654e-9
+ sky130_fd_pr__pfet_01v8__ua_diff_37 = -1.0238e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_37 = 0.27501
+ sky130_fd_pr__pfet_01v8__ub_diff_37 = 5.9384e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_37 = -0.0067074
+ sky130_fd_pr__pfet_01v8__pdits_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_37 = -0.11569
+ sky130_fd_pr__pfet_01v8__eta0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_37 = 0.0032138
+ sky130_fd_pr__pfet_01v8__vsat_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_37 = 0.020538
+ sky130_fd_pr__pfet_01v8__cgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_37 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 038, W = 0.42u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_38 = -7.3329e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_38 = 2.0396e-10
+ sky130_fd_pr__pfet_01v8__ua_diff_38 = -8.9609e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_38 = 0.27791
+ sky130_fd_pr__pfet_01v8__tvoff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_38 = 5.0883e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_38 = -0.012119
+ sky130_fd_pr__pfet_01v8__pdits_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_38 = -0.11437
+ sky130_fd_pr__pfet_01v8__eta0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_38 = 0.0029684
+ sky130_fd_pr__pfet_01v8__vsat_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_38 = -0.0074938
+ sky130_fd_pr__pfet_01v8__cgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_38 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 039, W = 0.42u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_39 = 1.0227e-7
+ sky130_fd_pr__pfet_01v8__agidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_39 = -4.0914e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_39 = -0.3
+ sky130_fd_pr__pfet_01v8__ua_diff_39 = -1.1205e-11
+ sky130_fd_pr__pfet_01v8__tvoff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_39 = -2.7333e-20
+ sky130_fd_pr__pfet_01v8__k2_diff_39 = 0.0074497
+ sky130_fd_pr__pfet_01v8__pdits_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_39 = -0.059118
+ sky130_fd_pr__pfet_01v8__eta0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_39 = 8.486e-5
+ sky130_fd_pr__pfet_01v8__vsat_diff_39 = 20005.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_39 = 0.049573
+ sky130_fd_pr__pfet_01v8__cgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_39 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 040, W = 0.42u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_40 = 1.348e-7
+ sky130_fd_pr__pfet_01v8__b1_diff_40 = 6.0708e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_40 = -4.4959e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_40 = 3.0442
+ sky130_fd_pr__pfet_01v8__ub_diff_40 = 4.1781e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_40 = -0.01793
+ sky130_fd_pr__pfet_01v8__voff_diff_40 = -0.17479
+ sky130_fd_pr__pfet_01v8__a0_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_40 = 18363.0
+ sky130_fd_pr__pfet_01v8__u0_diff_40 = 0.00070937
+ sky130_fd_pr__pfet_01v8__vth0_diff_40 = 0.020271
+ sky130_fd_pr__pfet_01v8__cgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_40 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 041, W = 0.42u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_41 = 5.5103e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_41 = 1.3639e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_41 = -4.6228e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_41 = 2.9421
+ sky130_fd_pr__pfet_01v8__ub_diff_41 = 4.5805e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_41 = -0.012839
+ sky130_fd_pr__pfet_01v8__voff_diff_41 = -0.26704
+ sky130_fd_pr__pfet_01v8__a0_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_41 = 19408.0
+ sky130_fd_pr__pfet_01v8__u0_diff_41 = 0.00082359
+ sky130_fd_pr__pfet_01v8__vth0_diff_41 = 0.049828
*
* sky130_fd_pr__pfet_01v8, Bin 042, W = 0.42u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__u0_diff_42 = 0.0019261
+ sky130_fd_pr__pfet_01v8__vth0_diff_42 = 0.02147
+ sky130_fd_pr__pfet_01v8__cgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_42 = -1.2525e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_42 = 4.1893e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_42 = -1.0522e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_42 = 0.57836
+ sky130_fd_pr__pfet_01v8__ub_diff_42 = 4.5194e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_42 = -0.0071804
+ sky130_fd_pr__pfet_01v8__voff_diff_42 = -0.17603
+ sky130_fd_pr__pfet_01v8__a0_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_42 = 20068.0
*
* sky130_fd_pr__pfet_01v8, Bin 043, W = 0.55u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_43 = 20090.0
+ sky130_fd_pr__pfet_01v8__u0_diff_43 = 0.0020132
+ sky130_fd_pr__pfet_01v8__vth0_diff_43 = -0.015677
+ sky130_fd_pr__pfet_01v8__cgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_43 = -2.0877e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_43 = -4.449e-10
+ sky130_fd_pr__pfet_01v8__agidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_43 = -1.0545e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_43 = 0.48051
+ sky130_fd_pr__pfet_01v8__ub_diff_43 = 3.9827e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_43 = -0.012381
+ sky130_fd_pr__pfet_01v8__voff_diff_43 = -0.13176
+ sky130_fd_pr__pfet_01v8__a0_diff_43 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 044, W = 0.55u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_44 = -0.10035
+ sky130_fd_pr__pfet_01v8__a0_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_44 = 0.0030032
+ sky130_fd_pr__pfet_01v8__vth0_diff_44 = 0.019075
+ sky130_fd_pr__pfet_01v8__cgidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_44 = -6.0544e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_44 = 4.9725e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_44 = 2.035e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_44 = 0.20225
+ sky130_fd_pr__pfet_01v8__ub_diff_44 = 5.5406e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_44 = -0.0089871
*
* sky130_fd_pr__pfet_01v8, Bin 045, W = 0.55u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_45 = 0.00042447
+ sky130_fd_pr__pfet_01v8__voff_diff_45 = -0.059301
+ sky130_fd_pr__pfet_01v8__a0_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_45 = 20022.0
+ sky130_fd_pr__pfet_01v8__u0_diff_45 = -0.00019504
+ sky130_fd_pr__pfet_01v8__vth0_diff_45 = 0.033581
+ sky130_fd_pr__pfet_01v8__cgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_45 = 8.8077e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_45 = 2.7625e-10
+ sky130_fd_pr__pfet_01v8__agidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_45 = -9.3232e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_45 = -0.1220159
+ sky130_fd_pr__pfet_01v8__ub_diff_45 = -3.8525e-20
*
* sky130_fd_pr__pfet_01v8, Bin 046, W = 0.55u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_46 = 0.4036
+ sky130_fd_pr__pfet_01v8__ub_diff_46 = 5.6923e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_46 = -0.013043
+ sky130_fd_pr__pfet_01v8__voff_diff_46 = -0.12363
+ sky130_fd_pr__pfet_01v8__a0_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_46 = 0.0033005
+ sky130_fd_pr__pfet_01v8__vsat_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_46 = -0.0040396
+ sky130_fd_pr__pfet_01v8__cgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_46 = -6.114e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_46 = 4.1551e-10
+ sky130_fd_pr__pfet_01v8__agidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_46 = -5.7212e-12
*
* sky130_fd_pr__pfet_01v8, Bin 047, W = 0.55u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_47 = 1.0557e-8
+ sky130_fd_pr__pfet_01v8__ua_diff_47 = -4.5957e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_47 = 2.7386
+ sky130_fd_pr__pfet_01v8__ub_diff_47 = 4.3457e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_47 = -0.0056125
+ sky130_fd_pr__pfet_01v8__voff_diff_47 = -0.22548
+ sky130_fd_pr__pfet_01v8__eta0_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_47 = 0.00069904
+ sky130_fd_pr__pfet_01v8__vsat_diff_47 = 19768.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_47 = 0.006925
+ sky130_fd_pr__pfet_01v8__cgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_47 = 3.8587e-7
*
* sky130_fd_pr__pfet_01v8, Bin 048, W = 0.55u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_48 = -3.1638e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_48 = -5.283e-10
+ sky130_fd_pr__pfet_01v8__ua_diff_48 = -7.9455e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_48 = 0.27288
+ sky130_fd_pr__pfet_01v8__ub_diff_48 = 4.129e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_48 = -0.017392
+ sky130_fd_pr__pfet_01v8__pdits_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_48 = -0.13858
+ sky130_fd_pr__pfet_01v8__eta0_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_48 = 0.0016268
+ sky130_fd_pr__pfet_01v8__vsat_diff_48 = 20057.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_48 = 0.026387
+ sky130_fd_pr__pfet_01v8__cgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_48 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 049, W = 0.64u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_49 = 4.7891e-7
+ sky130_fd_pr__pfet_01v8__agidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_49 = 2.8741e-9
+ sky130_fd_pr__pfet_01v8__ua_diff_49 = -1.5419e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_49 = 3.2565
+ sky130_fd_pr__pfet_01v8__tvoff_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_49 = 4.4353e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_49 = -0.00076033
+ sky130_fd_pr__pfet_01v8__pdits_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_49 = -0.042312
+ sky130_fd_pr__pfet_01v8__eta0_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_49 = 0.00030997
+ sky130_fd_pr__pfet_01v8__vsat_diff_49 = 22556.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_49 = -0.083901
+ sky130_fd_pr__pfet_01v8__cgidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_49 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 050, W = 0.84u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_50 = -1.2127e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_50 = 2.6465
+ sky130_fd_pr__pfet_01v8__ub_diff_50 = 4.4559e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_50 = -0.033534
+ sky130_fd_pr__pfet_01v8__voff_diff_50 = -0.13229
+ sky130_fd_pr__pfet_01v8__a0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_50 = -10846.0
+ sky130_fd_pr__pfet_01v8__u0_diff_50 = 0.00055104
+ sky130_fd_pr__pfet_01v8__vth0_diff_50 = -0.092463
+ sky130_fd_pr__pfet_01v8__cgidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_50 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 051, W = 1.65u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_51 = -4.2859e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_51 = 2.0274
+ sky130_fd_pr__pfet_01v8__ub_diff_51 = 2.55e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_51 = -0.014919
+ sky130_fd_pr__pfet_01v8__voff_diff_51 = -0.18661
+ sky130_fd_pr__pfet_01v8__a0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_51 = -7007.1
+ sky130_fd_pr__pfet_01v8__u0_diff_51 = 0.00037115
+ sky130_fd_pr__pfet_01v8__vth0_diff_51 = -0.060745
+ sky130_fd_pr__pfet_01v8__cgidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_51 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8.pm3.spice"
