* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 38
.param
+ sky130_fd_pr__nfet_01v8_lvt__toxe_mult = 1.0
+ sky130_fd_pr__nfet_01v8_lvt__rshn_mult = 1.0
+ sky130_fd_pr__nfet_01v8_lvt__overlap_mult = 0.92429
+ sky130_fd_pr__nfet_01v8_lvt__ajunction_mult = 1.0004
+ sky130_fd_pr__nfet_01v8_lvt__pjunction_mult = 0.89176
+ sky130_fd_pr__nfet_01v8_lvt__lint_diff = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__wint_diff = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__dlc_diff = -1.3619e-9
+ sky130_fd_pr__nfet_01v8_lvt__dwc_diff = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 000, W = 1.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_0 = -0.061491
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_0 = -0.047706
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_0 = 0.0081568
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_0 = 0.00022078
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0 = 0.0018585
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_0 = -0.097377
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_0 = 6.4377e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_0 = 2.3269e-19
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0 = 0.20403
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0 = 0.00049577
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 001, W = 1.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_1 = -0.064357
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_1 = -0.048796
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_1 = 0.0073323
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1 = 0.001658
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_1 = -0.13298
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_1 = -0.00089095
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_1 = 3.5508e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_1 = 1.8212e-19
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1 = 0.20651
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1 = -0.0026634
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 002, W = 1.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2 = -0.00074866
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_2 = -0.0047222
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_2 = -0.066564
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_2 = 0.0097539
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2 = -0.0003155
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_2 = 0.028996
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_2 = -0.0011451
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_2 = -6.2443e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_2 = 1.6879e-19
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2 = 0.26551
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 003, W = 1.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3 = 0.33579
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3 = 0.025971
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_3 = -0.055736
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_3 = 0.0025471
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3 = -0.00014158
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_3 = 0.00072662
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_3 = -1.4438e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3 = -10.8
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_3 = 1.6748e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 004, W = 1.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4 = 0.43618
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4 = 0.0058944
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_4 = -0.070254
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_4 = 0.0019871
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4 = 0.00034993
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_4 = -0.00078107
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_4 = 2.7231e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4 = 1469.3
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_4 = 4.4948e-22
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 005, W = 1.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_5 = 1.8383e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5 = 0.39129
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5 = 0.019258
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_5 = -0.073895
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_5 = 0.0054573
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5 = 0.0011151
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_5 = -0.00049991
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_5 = -1.444e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5 = -5412.1
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_5 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 006, W = 1.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_6 = 1.2732e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6 = 0.26849
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6 = 0.00059786
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_6 = -0.055874
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_6 = 0.001201
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6 = 0.0018628
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_6 = -0.00033778
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_6 = -5.5154e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6 = 5238.9
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_6 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 007, W = 3.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_7 = 1.5266e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7 = 0.13341
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7 = 0.0046366
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_7 = -0.047492
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_7 = -0.030992
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_7 = 0.0048651
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7 = 0.0023604
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_7 = -0.054999
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_7 = 0.0007892
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_7 = -1.2977e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 008, W = 3.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8 = 0.0028337
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_8 = -0.07263
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_8 = 0.00056632
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_8 = 4.2479e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_8 = 1.7315e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8 = 0.13375
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8 = -0.0037694
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_8 = -0.049464
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_8 = -0.032894
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_8 = 0.0029323
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 009, W = 3.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9 = 0.0025089
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_9 = -0.0069325
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_9 = -6.5502e-5
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_9 = -9.0975e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_9 = 1.0671e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9 = 0.16029
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9 = 3.5662e-5
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_9 = 0.001561
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_9 = -0.038551
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_9 = 0.0064203
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 010, W = 3.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_10 = 3.9245e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_10 = -3.2886e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10 = 0.001867
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_10 = -0.0014665
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10 = 3984.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10 = -0.012631
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10 = -0.033459
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_10 = -0.0028083
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_10 = 0.003079
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 011, W = 3.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_11 = 0.0042111
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_11 = 1.1147e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_11 = 1.6097e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11 = -0.00088129
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_11 = 0.0010862
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11 = 7628.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11 = 0.010789
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11 = 0.46349
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_11 = -0.065727
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 012, W = 3.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_12 = 0.0077253
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_12 = 1.6468e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_12 = 2.4517e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12 = -0.00028352
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_12 = 0.00015296
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12 = 5086.2
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12 = 0.010933
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12 = 0.35367
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_12 = -0.063364
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_12 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 013, W = 3.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_13 = 0.01115
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_13 = -1.213e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_13 = 1.8252e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13 = 0.0024997
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_13 = 0.00086105
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13 = 9243.7
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13 = 0.0081041
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13 = 0.2278
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_13 = -0.038891
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_13 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 014, W = 5.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14 = 0.071645
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_14 = -0.023211
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_14 = 0.0032333
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_14 = -6.8844e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_14 = 1.7832e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_14 = -0.054744
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14 = 0.003378
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_14 = -0.073674
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_14 = 0.001075
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14 = -0.0032136
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 015, W = 5.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15 = 0.0033883
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15 = 0.14879
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_15 = -0.031961
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_15 = -0.0058846
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_15 = -1.4976e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_15 = 1.8105e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_15 = -0.0057138
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15 = 0.0026718
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_15 = -0.015857
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_15 = 0.00082745
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 016, W = 5.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16 = 0.0027459
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_16 = -0.045808
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_16 = 0.00041893
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16 = -0.0070266
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16 = 0.10789
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_16 = -0.025262
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_16 = 0.009614
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_16 = 1.8675e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_16 = 1.4212e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_16 = 0.0059522
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 017, W = 5.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17 = 0.0040963
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_17 = 0.00091908
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17 = 7738.8
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17 = -0.0056655
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17 = 0.19202
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_17 = -0.026515
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_17 = 0.002832
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_17 = -1.0056e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_17 = 1.9308e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 018, W = 5.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18 = 0.0024469
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_18 = 0.00014169
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18 = 1320.7
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18 = 0.01696
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18 = 0.28978
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_18 = -0.023719
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_18 = 0.0049699
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_18 = 1.6514e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_18 = 1.2088e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 019, W = 5.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_19 = 1.6091e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19 = 0.0024504
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_19 = -0.0013187
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19 = -2131.7
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19 = -0.0011996
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19 = 0.23158
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_19 = -0.040948
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_19 = 0.0054353
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_19 = 3.4787e-12
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 020, W = 5.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_20 = -3.3561e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_20 = 2.4427e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20 = 0.0030468
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_20 = 0.001822
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20 = 10521.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20 = -0.0006357
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20 = 0.19214
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_20 = -0.029574
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_20 = 0.0030478
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 021, W = 7.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_21 = -2.7372e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_21 = 2.0476e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_21 = 0.0069635
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21 = 0.0021399
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_21 = 0.0079875
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_21 = 0.0014395
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21 = 0.0052151
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21 = 0.17006
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_21 = -0.03417
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_21 = -0.0035982
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 022, W = 7.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_22 = 0.0085737
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_22 = -7.0145e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_22 = 1.5875e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_22 = -0.024942
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22 = 0.003229
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_22 = -0.056733
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_22 = 0.00072081
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22 = -0.0023361
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22 = 0.10855
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_22 = -0.024398
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 023, W = 7.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_23 = 0.007571
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_23 = -2.3602e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_23 = 2.0151e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_23 = -0.00081114
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23 = 0.00056944
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_23 = 0.01152
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_23 = 0.0009344
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23 = -0.0023254
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23 = 0.1891
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_23 = -0.04963
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_23 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 024, W = 7.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_24 = 0.0085689
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_24 = 6.3921e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_24 = -1.368e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24 = 0.0045
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_24 = -0.0026537
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24 = 6227.6
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24 = -0.01413
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24 = -0.0076286
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_24 = -0.0049977
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_24 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 025, W = 7.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25 = 0.31419
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_25 = -0.021009
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_25 = 0.006586
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_25 = 2.7798e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_25 = 1.0889e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25 = 0.0039624
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_25 = 7.4777e-5
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25 = 5048.1
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25 = 0.0065429
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 026, W = 7.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26 = 0.0018791
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26 = 0.23224
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_26 = -0.035392
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_26 = 0.0067513
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_26 = 1.7984e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_26 = 2.6984e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26 = 0.0026663
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_26 = -9.2827e-5
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26 = 4536.6
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 027, W = 7.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27 = 0.0031138
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_27 = 0.001424
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27 = 887.27
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27 = 0.0045997
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27 = 0.16118
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_27 = -0.026893
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_27 = 0.0039291
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_27 = -3.9545e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_27 = 2.1162e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 028, W = 0.42u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28 = 0.0014482
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_28 = -0.0019991
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28 = -0.0072946
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28 = 0.22299
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_28 = -0.052006
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_28 = 7.6327e-8
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_28 = 2.6382e-9
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_28 = 0.00271
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_28 = 2.8232e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_28 = 2.5216e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 029, W = 0.42u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29 = 0.00072929
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_29 = 0.00019904
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29 = 12088.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29 = 0.028839
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29 = 0.65782
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_29 = -0.090911
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_29 = 0.0010093
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_29 = 7.1505e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_29 = -3.5996e-20
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 030, W = 0.42u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_30 = 4.6407e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30 = -0.00024137
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_30 = 0.00097317
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30 = -166.39
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30 = -0.028905
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30 = 0.43815
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_30 = -0.080495
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_30 = -0.00080889
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_30 = 4.4458e-12
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 031, W = 0.55u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_31 = 1.5736e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_31 = -2.585e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31 = -0.00024285
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_31 = -0.00082845
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31 = 3589.6
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31 = 0.03604
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31 = 0.65757
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_31 = -0.090978
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_31 = -0.0031204
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 032, W = 0.64u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_32 = 1.2811e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_32 = -1.4693e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32 = -0.00081158
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_32 = -0.00032917
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32 = 10009.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32 = 0.025783
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32 = 0.58301
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_32 = -0.070773
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_32 = -0.0040461
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 033, W = 0.84u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_33 = -0.0049622
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_33 = 8.2057e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_33 = -1.3909e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33 = -0.00029263
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_33 = -0.00039887
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33 = 10623.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33 = 0.03326
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33 = 0.65685
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_33 = -0.080184
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 034, W = 1.65u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_34 = 0.030843
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_34 = 6.5406e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_34 = -2.2057e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34 = -0.00088378
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_34 = -0.0020042
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34 = 6655.9
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34 = 0.0053876
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34 = 0.30472
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_34 = -0.015046
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_34 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 035, W = 3.01u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_35 = 0.023992
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_35 = 4.3469e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_35 = -1.4528e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35 = -0.00075682
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_35 = -0.0016712
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35 = 3027.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35 = -0.0028534
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35 = 0.1846
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_35 = -0.018025
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_35 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 036, W = 5.05u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36 = 0.2588
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_36 = -0.043593
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_36 = 0.025521
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_36 = 1.3825e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_36 = 5.9588e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36 = 0.0021024
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_36 = -0.00039882
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36 = 8556.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36 = -0.0026425
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 037, W = 5.05u, L = 0.25u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37 = -6.3651e-5
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37 = 0.24722
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_37 = -0.044109
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_37 = 0.019583
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_37 = 2.1451e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_37 = -1.4683e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37 = 0.002514
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_37 = -0.0040277
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37 = 172.72
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_01v8_lvt.pm3.spice"
