* SKY130 Spice File.
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_01v8__tt.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_01v8_lvt__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8_lvt__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_g5v0d10v5__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_g5v0d10v5__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice"
.include "sky130_fd_pr_models/corners/tt/nonfet.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_20v0__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_20v0__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_20v0_nvt__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/all.spice"
.include "sky130_fd_pr_models/corners/tt/rf.spice"
