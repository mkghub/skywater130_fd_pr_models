* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff = -0.0850
* Number of bins: 40
.param
+ sky130_fd_pr__pfet_01v8_lvt__toxe_mult = 1.0
+ sky130_fd_pr__pfet_01v8_lvt__rshp_mult = 1.0
+ sky130_fd_pr__pfet_01v8_lvt__overlap_mult = 0.2
+ sky130_fd_pr__pfet_01v8_lvt__ajunction_mult = 9.9626e-1
+ sky130_fd_pr__pfet_01v8_lvt__pjunction_mult = 1.0009e+0
+ sky130_fd_pr__pfet_01v8_lvt__lint_diff = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__wint_diff = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__dlc_diff = -12.0e-9
+ sky130_fd_pr__pfet_01v8_lvt__dwc_diff = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 000, W = 1.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_0 = 2.1451e-5
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_0 = 0.17464
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_0 = ' -0.045471 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_0 = 0.060517
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_0 = 0.0071015
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 001, W = 1.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_1 = -0.00030403
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_1 = 2.0909e-5
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_1 = 0.12938
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_1 = ' -0.013221 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_1 = 0.089162
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 002, W = 1.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_2 = 0.11464
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_2 = 0.0045081
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_2 = -7.5619e-5
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_2 = 0.067503
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_2 = ' -0.0096086 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_2 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 003, W = 1.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_3 = 0.093146
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_3 = -0.0012403
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_3 = 1.7182e-5
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_3 = 0.11591
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_3 = ' -0.023987 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 004, W = 1.0u, L = 0.35u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_4 = ' -0.093844 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_4 = -1.7546e-7
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_4 = -0.011657
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_4 = -7.0716e-5
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_4 = 16031.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_4 = 2.0585e-7
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_4 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 005, W = 1.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_5 = ' -0.023527 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_5 = -1.102e-7
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_5 = -0.0044621
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_5 = -2.4829e-5
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_5 = -19187.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_5 = 1.1181e-7
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_5 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 006, W = 3.0u, L = 1.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_6 = 0.26426
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_6 = ' -0.04313 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_6 = 0.01788
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_6 = -0.0019941
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_6 = -0.00016957
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_6 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 007, W = 3.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_7 = 0.23041
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_7 = ' -0.041229 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_7 = 0.064964
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_7 = 0.0011069
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_7 = -1.4444e-5
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_7 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 008, W = 3.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_8 = 0.20351
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_8 = ' -0.014884 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_8 = 0.053383
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_8 = 0.001511
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_8 = -0.00019792
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_8 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 009, W = 3.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_9 = 0.18803
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_9 = ' -0.021303 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_9 = 0.073088
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_9 = 0.0054858
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_9 = -0.00019305
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_9 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 010, W = 3.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_10 = -0.00015805
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_10 = ' -0.0097702 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_10 = 0.0014514
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_10 = 0.11926
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_10 = 0.094176
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 011, W = 3.0u, L = 0.35u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_11 = -0.00019399
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_11 = 18916.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_11 = ' -0.047588 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_11 = 0.0078636
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_11 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 012, W = 3.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_12 = -0.00046191
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_12 = 0.077339
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_12 = -0.000237
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_12 = -6368.4
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_12 = ' -0.029472 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_12 = -1.0985e-6
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_12 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 013, W = 5.0u, L = 1.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_13 = -0.0002228
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_13 = 0.085125
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_13 = 0.10287
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_13 = -8.1063e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_13 = ' -0.024537 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_13 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 014, W = 5.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_14 = 0.00021102
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_14 = 0.078811
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_14 = 0.1086
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_14 = 9.4292e-6
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_14 = ' -0.032734 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_14 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 015, W = 5.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_15 = 0.0012137
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_15 = 0.10136
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_15 = 0.10469
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_15 = -6.6693e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_15 = ' -0.028044 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_15 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 016, W = 5.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_16 = 0.0019673
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_16 = 0.083685
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_16 = 0.10692
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_16 = -7.4938e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_16 = ' -0.020294 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_16 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 017, W = 5.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_17 = 0.0025126
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_17 = 0.094989
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_17 = 0.10267
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_17 = -9.6003e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_17 = ' -0.01386 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_17 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 018, W = 5.0u, L = 0.35u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_18 = 0.0035857
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_18 = -7.1375e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_18 = 8295.2
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_18 = ' -0.066303 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_18 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 019, W = 5.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_19 = -1.2407e-6
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_19 = -0.0036875
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_19 = 0.058101
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_19 = -2.1001e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_19 = -9997.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_19 = ' -0.057784 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 020, W = 7.0u, L = 1.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_20 = -0.0074997
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_20 = 0.18147
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_20 = 0.047551
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_20 = -2.3889e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_20 = ' -0.043041 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 021, W = 7.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_21 = -2.3186e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_21 = ' -0.044365 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_21 = -0.0033081
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_21 = 0.21309
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_21 = 0.073049
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 022, W = 7.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_22 = 0.21951
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_22 = 0.060844
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_22 = 7.3356e-6
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_22 = ' -0.045242 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__uc_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_22 = -0.0054151
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_22 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 023, W = 7.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_23 = 0.0016295
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_23 = 0.049924
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_23 = 0.11673
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_23 = -1.8122e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_23 = ' -0.023069 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_23 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 024, W = 7.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_24 = 0.00051387
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_24 = 0.068356
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_24 = 0.11339
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_24 = 8.2839e-6
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_24 = ' -0.032509 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_24 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 025, W = 7.0u, L = 0.35u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_25 = 0.0014271
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_25 = 1.3336e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_25 = 10704.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_25 = ' -0.079917 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_25 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 026, W = 7.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_26 = -0.0044363
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_26 = 0.067715
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_26 = -4.0559e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_26 = 12124.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_26 = ' -0.045124 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_26 = -7.3883e-7
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 027, W = 0.42u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_27 = -1.6046e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_27 = 4.4049e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_27 = -0.0079686
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_27 = 0.00048641
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_27 = ' -0.094912 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_27 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 028, W = 0.42u, L = 20.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_28 = -1.3014e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_28 = 2.2895e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_28 = -0.0062032
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_28 = -7.101e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_28 = ' -0.0027948 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_28 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 029, W = 0.42u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_29 = -1.1083e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_29 = 2.2784e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_29 = -0.0071632
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_29 = 1.223e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_29 = ' -0.013234 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_29 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 030, W = 0.42u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_30 = -1.226e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_30 = 2.4821e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_30 = -0.0055578
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_30 = 6.2391e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_30 = ' -0.032311 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_30 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 031, W = 0.42u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_31 = -5.34e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_31 = 2.2699e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_31 = -0.0037977
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_31 = -3.489e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_31 = ' -0.0014815 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 032, W = 0.42u, L = 0.35u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_32 = 2.7696e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_32 = 15069.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_32 = ' 0.029512 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_32 = 0.0080418
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_32 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 033, W = 0.42u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_33 = 4.0289e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_33 = -17161.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_33 = ' -0.058342 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_33 = -1.8961e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_33 = 2.1168e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_33 = -0.012786
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_33 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 034, W = 0.55u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_34 = 0.0016548
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_34 = 3.3603e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_34 = ' -0.0087662 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_34 = -7.52e-8
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_34 = 3.435e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_34 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 035, W = 0.55u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_35 = 0.011772
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_35 = 3.5846e-5
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_35 = ' -0.02365 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_35 = -1.0503e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_35 = 2.0297e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_35 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 036, W = 0.55u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_36 = 0.011867
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_36 = 1.6269e-6
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_36 = ' -0.026415 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_36 = -1.4822e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_36 = 2.0228e-7
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 037, W = 0.55u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_37 = 2.0418e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_37 = 0.0090638
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_37 = -6.574e-6
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_37 = ' -0.018088 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_37 = -8.3896e-8
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 038, W = 0.55u, L = 0.35u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_38 = -0.0055494
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_38 = 0.00010812
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_38 = 17194.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_38 = ' -0.10569 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_38 = 0.0
*
* sky130_fd_pr__pfet_01v8_lvt, Bin 039, W = 0.55u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8_lvt__pclm_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kt1_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b0_diff_39 = -1.7931e-7
+ sky130_fd_pr__pfet_01v8_lvt__pdits_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__b1_diff_39 = 4.118e-7
+ sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__agidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ub_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__voff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__k2_diff_39 = -0.019137
+ sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__eta0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ags_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__a0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__u0_diff_39 = 0.00035271
+ sky130_fd_pr__pfet_01v8_lvt__vsat_diff_39 = -15626.0
+ sky130_fd_pr__pfet_01v8_lvt__vth0_diff_39 = ' -0.12364 + sky130_fd_pr__pfet_01v8_lvt__vth0_correldiff'
+ sky130_fd_pr__pfet_01v8_lvt__keta_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__ua_diff_39 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8_lvt.pm3.spice"
