* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 11
.param
+ sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult = 0.958
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult = 1.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult = 0.80232
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult = 8.7078e-1
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult = 8.4883e-1
+ sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff = 1.21275e-8
+ sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff = -2.252e-8
+ sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff = 1.21275e-8
+ sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff = -2.252e-8
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 000, W = 17.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_0 = 0.16357
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_0 = 0.0029504
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_0 = 0.00101
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_0 = 0.0011108
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_0 = -4523.2
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_0 = -7.1223e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_0 = -2.3306e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_0 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_0 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 001, W = 19.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_1 = 0.17171
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_1 = 0.0035138
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_1 = 0.0027963
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_1 = 0.0025467
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_1 = -4339.5
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_1 = -6.2712e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_1 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_1 = -3.9765e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_1 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 002, W = 21.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_2 = 0.17982
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_2 = 0.0032498
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_2 = 0.0011356
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_2 = 0.0016785
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_2 = -2873.5
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_2 = -6.3605e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_2 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_2 = -1.631e-11
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 003, W = 23.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_3 = -1.1281e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_3 = 0.17002
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_3 = 0.0032597
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_3 = 0.0009255
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_3 = 0.002901
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_3 = -2782.4
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_3 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_3 = -6.483e-19
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 004, W = 26.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_4 = -6.9589e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_4 = -2.3104e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_4 = 0.16286
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_4 = 0.0012986
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_4 = 0.0012232
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_4 = 0.00053733
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_4 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_4 = -3682.5
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_4 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 005, W = 30.25u, L = 1.0u
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_5 = -9.6362e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_5 = 1.0425e-10
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_5 = 0.19678
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_5 = 0.1098
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_5 = -0.4
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_5 = 0.051952
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_5 = -0.0049958
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_5 = 0.0039808
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_5 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_5 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 006, W = 30.25u, L = 0.55u
* ------------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_6 = -3.9259e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_6 = -2.2649e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_6 = 0.16025
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_6 = 0.0023857
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_6 = 0.00149
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_6 = 0.00087375
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_6 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_6 = -1484.1
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 007, W = 40.31u, L = 0.55u
* ------------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_7 = -116.16
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_7 = -6.7577e-20
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_7 = -6.9305e-12
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_7 = 0.13958
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_7 = 0.002226
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_7 = 0.0012851
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_7 = 0.0021027
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 008, W = 50.99u, L = 1.0u
* -----------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_8 = -0.0075657
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_8 = 0.00029955
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_8 = -1.1175e-18
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_8 = 9.2607e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_8 = 0.19208
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_8 = 0.07794
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_8 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_8 = -0.3401
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_8 = 0.014154
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 009, W = 50.99u, L = 0.55u
* ------------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_9 = -0.0036012
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_9 = 0.0035682
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_9 = -0.0063521
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_9 = -3184.4
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_9 = 2.4123e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_9 = -3.0465e-11
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_9 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_9 = 0.14429
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_9 = 0.0
*
* sky130_fd_pr__esd_nfet_g5v0d10v5, Bin 010, W = 5.4u, L = 0.6u
* ---------------------------------
+ sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_10 = -1.2342e-12
+ sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_10 = -4918.4
+ sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_10 = -4.9751e-19
+ sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_10 = -0.0011713
+ sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_10 = 0.27905
+ sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_10 = -0.00098474
+ sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_10 = 0.00297
+ sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_10 = 0.0
+ sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_10 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice"
