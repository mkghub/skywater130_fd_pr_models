* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 63
.param
+ sky130_fd_pr__nfet_01v8__toxe_mult = 1.0365
+ sky130_fd_pr__nfet_01v8__rshn_mult = 1.0
+ sky130_fd_pr__nfet_01v8__overlap_mult = 0.98
+ sky130_fd_pr__nfet_01v8__lint_diff = -1.21275e-8
+ sky130_fd_pr__nfet_01v8__wint_diff = 2.252e-8
+ sky130_fd_pr__nfet_01v8__dlc_diff = -11.107e-9
+ sky130_fd_pr__nfet_01v8__dwc_diff = 2.252e-8
*
* sky130_fd_pr__nfet_01v8, Bin 000, W = 1.26u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__voff_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_0 = -1.549e-19
+ sky130_fd_pr__nfet_01v8__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_0 = 3.6167e-11
+ sky130_fd_pr__nfet_01v8__vsat_diff_0 = 34157.0
+ sky130_fd_pr__nfet_01v8__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_0 = -0.017901
+ sky130_fd_pr__nfet_01v8__vth0_diff_0 = 0.030223
+ sky130_fd_pr__nfet_01v8__nfactor_diff_0 = -0.0030628
+ sky130_fd_pr__nfet_01v8__u0_diff_0 = -0.0026696
+ sky130_fd_pr__nfet_01v8__eta0_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_0 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 001, W = 1.68u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_1 = -3.8533e-19
+ sky130_fd_pr__nfet_01v8__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_1 = 1.055e-10
+ sky130_fd_pr__nfet_01v8__vsat_diff_1 = 15769.0
+ sky130_fd_pr__nfet_01v8__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_1 = -0.013558
+ sky130_fd_pr__nfet_01v8__vth0_diff_1 = 0.06096
+ sky130_fd_pr__nfet_01v8__nfactor_diff_1 = -0.18837
+ sky130_fd_pr__nfet_01v8__u0_diff_1 = -0.0015015
*
* sky130_fd_pr__nfet_01v8, Bin 002, W = 1.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__nfactor_diff_2 = 1.0676
+ sky130_fd_pr__nfet_01v8__u0_diff_2 = -0.0023051
+ sky130_fd_pr__nfet_01v8__vth0_diff_2 = 0.013135
+ sky130_fd_pr__nfet_01v8__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_2 = 5.2609e-21
+ sky130_fd_pr__nfet_01v8__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_2 = 7.974e-12
+ sky130_fd_pr__nfet_01v8__vsat_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_2 = -0.054816
+ sky130_fd_pr__nfet_01v8__a0_diff_2 = 0.2494
+ sky130_fd_pr__nfet_01v8__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_2 = -0.0074533
*
* sky130_fd_pr__nfet_01v8, Bin 003, W = 1.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_3 = -0.0057524
+ sky130_fd_pr__nfet_01v8__nfactor_diff_3 = 0.78012
+ sky130_fd_pr__nfet_01v8__u0_diff_3 = -0.0022191
+ sky130_fd_pr__nfet_01v8__vth0_diff_3 = 0.0042677
+ sky130_fd_pr__nfet_01v8__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_3 = -9.5237e-20
+ sky130_fd_pr__nfet_01v8__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_3 = 5.8568e-12
+ sky130_fd_pr__nfet_01v8__vsat_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_3 = -0.0010882
+ sky130_fd_pr__nfet_01v8__a0_diff_3 = 0.020299
+ sky130_fd_pr__nfet_01v8__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_3 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 004, W = 1.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_4 = 0.0048793
+ sky130_fd_pr__nfet_01v8__nfactor_diff_4 = 1.1419
+ sky130_fd_pr__nfet_01v8__u0_diff_4 = -0.0029667
+ sky130_fd_pr__nfet_01v8__vth0_diff_4 = -0.0051998
+ sky130_fd_pr__nfet_01v8__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_4 = -1.7579e-19
+ sky130_fd_pr__nfet_01v8__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_4 = 6.8705e-12
+ sky130_fd_pr__nfet_01v8__vsat_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_4 = -0.026541
+ sky130_fd_pr__nfet_01v8__a0_diff_4 = 0.069075
+ sky130_fd_pr__nfet_01v8__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_4 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 005, W = 1.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_5 = 0.0075232
+ sky130_fd_pr__nfet_01v8__nfactor_diff_5 = 1.3493
+ sky130_fd_pr__nfet_01v8__u0_diff_5 = -0.0035065
+ sky130_fd_pr__nfet_01v8__vth0_diff_5 = -0.010021
+ sky130_fd_pr__nfet_01v8__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_5 = -1.8081e-19
+ sky130_fd_pr__nfet_01v8__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_5 = 8.4463e-12
+ sky130_fd_pr__nfet_01v8__vsat_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_5 = -0.029492
+ sky130_fd_pr__nfet_01v8__a0_diff_5 = 0.068611
+ sky130_fd_pr__nfet_01v8__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_5 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 006, W = 1.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_6 = -0.020268
+ sky130_fd_pr__nfet_01v8__nfactor_diff_6 = 0.39175
+ sky130_fd_pr__nfet_01v8__u0_diff_6 = -0.0031675
+ sky130_fd_pr__nfet_01v8__vth0_diff_6 = 0.055773
+ sky130_fd_pr__nfet_01v8__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_6 = -6.466e-19
+ sky130_fd_pr__nfet_01v8__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_6 = 1.1729e-10
+ sky130_fd_pr__nfet_01v8__vsat_diff_6 = 21852.0
+ sky130_fd_pr__nfet_01v8__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_6 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 007, W = 1.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_7 = -0.010135
+ sky130_fd_pr__nfet_01v8__nfactor_diff_7 = -0.37696
+ sky130_fd_pr__nfet_01v8__u0_diff_7 = -0.0052365
+ sky130_fd_pr__nfet_01v8__vth0_diff_7 = 0.0259
+ sky130_fd_pr__nfet_01v8__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_7 = -6.349e-19
+ sky130_fd_pr__nfet_01v8__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_7 = 1.0396e-10
+ sky130_fd_pr__nfet_01v8__vsat_diff_7 = 22273.0
+ sky130_fd_pr__nfet_01v8__a0_diff_7 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 008, W = 1.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__a0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_8 = 8.156e-11
+ sky130_fd_pr__nfet_01v8__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_8 = -0.0051255
+ sky130_fd_pr__nfet_01v8__nfactor_diff_8 = 0.73062
+ sky130_fd_pr__nfet_01v8__u0_diff_8 = -0.011342
+ sky130_fd_pr__nfet_01v8__vth0_diff_8 = 0.0082733
+ sky130_fd_pr__nfet_01v8__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_8 = -6.9309e-19
+ sky130_fd_pr__nfet_01v8__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_8 = 8930.1
*
* sky130_fd_pr__nfet_01v8, Bin 009, W = 1.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__kt1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_9 = -2.577e-19
+ sky130_fd_pr__nfet_01v8__vsat_diff_9 = 5776.5
+ sky130_fd_pr__nfet_01v8__a0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_9 = 9.8611e-12
+ sky130_fd_pr__nfet_01v8__tvoff_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_9 = 0.0042009
+ sky130_fd_pr__nfet_01v8__nfactor_diff_9 = 1.3748
+ sky130_fd_pr__nfet_01v8__u0_diff_9 = -0.0037139
+ sky130_fd_pr__nfet_01v8__vth0_diff_9 = 0.010066
+ sky130_fd_pr__nfet_01v8__eta0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_9 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 010, W = 2.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__ags_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_10 = -0.018067
+ sky130_fd_pr__nfet_01v8__ua_diff_10 = 7.6823e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_10 = -3.4649e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_10 = 16146.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_10 = 0.053513
+ sky130_fd_pr__nfet_01v8__pdits_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_10 = 0.27497
+ sky130_fd_pr__nfet_01v8__u0_diff_10 = -0.00026336
*
* sky130_fd_pr__nfet_01v8, Bin 011, W = 3.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__pclm_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_11 = 1.0158
+ sky130_fd_pr__nfet_01v8__u0_diff_11 = -0.0012241
+ sky130_fd_pr__nfet_01v8__ags_diff_11 = -0.055378
+ sky130_fd_pr__nfet_01v8__keta_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_11 = -0.0043261
+ sky130_fd_pr__nfet_01v8__ua_diff_11 = 3.2122e-12
+ sky130_fd_pr__nfet_01v8__eta0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_11 = -5.662e-20
+ sky130_fd_pr__nfet_01v8__tvoff_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_11 = 0.023173
+ sky130_fd_pr__nfet_01v8__rdsw_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_11 = 0.0080793
+ sky130_fd_pr__nfet_01v8__pdits_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_11 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 012, W = 3.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__pditsd_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_12 = 1.0006
+ sky130_fd_pr__nfet_01v8__u0_diff_12 = -0.0042244
+ sky130_fd_pr__nfet_01v8__ags_diff_12 = -0.091091
+ sky130_fd_pr__nfet_01v8__keta_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_12 = 0.003506
+ sky130_fd_pr__nfet_01v8__ua_diff_12 = 1.0697e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_12 = -4.0264e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_12 = 0.094702
+ sky130_fd_pr__nfet_01v8__rdsw_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_12 = -0.011754
+ sky130_fd_pr__nfet_01v8__pdits_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_12 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 013, W = 3.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__pdits_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_13 = 0.66116
+ sky130_fd_pr__nfet_01v8__u0_diff_13 = -0.0031486
+ sky130_fd_pr__nfet_01v8__ags_diff_13 = -0.042324
+ sky130_fd_pr__nfet_01v8__keta_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_13 = 0.0022844
+ sky130_fd_pr__nfet_01v8__ua_diff_13 = 1.5301e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_13 = -2.7829e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_13 = 0.07794
+ sky130_fd_pr__nfet_01v8__rdsw_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_13 = -0.0039027
+ sky130_fd_pr__nfet_01v8__b0_diff_13 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 014, W = 3.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__b0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_14 = 0.73725
+ sky130_fd_pr__nfet_01v8__u0_diff_14 = -0.0027435
+ sky130_fd_pr__nfet_01v8__ags_diff_14 = -0.057244
+ sky130_fd_pr__nfet_01v8__keta_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_14 = 0.0034323
+ sky130_fd_pr__nfet_01v8__ua_diff_14 = 6.7647e-12
+ sky130_fd_pr__nfet_01v8__eta0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_14 = -2.5224e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_14 = 0.080908
+ sky130_fd_pr__nfet_01v8__rdsw_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_14 = -0.0073519
*
* sky130_fd_pr__nfet_01v8, Bin 015, W = 3.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__kt1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_15 = 18445.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_15 = 0.028937
+ sky130_fd_pr__nfet_01v8__b0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_15 = 0.9748
+ sky130_fd_pr__nfet_01v8__u0_diff_15 = -0.0020123
+ sky130_fd_pr__nfet_01v8__ags_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_15 = -0.010671
+ sky130_fd_pr__nfet_01v8__ua_diff_15 = 1.2877e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_15 = -2.6848e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_15 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 016, W = 3.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__a0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_16 = 19149.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_16 = 0.024877
+ sky130_fd_pr__nfet_01v8__b0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_16 = 0.77183
+ sky130_fd_pr__nfet_01v8__u0_diff_16 = -0.0023051
+ sky130_fd_pr__nfet_01v8__ags_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_16 = -0.0062094
+ sky130_fd_pr__nfet_01v8__ua_diff_16 = 1.6209e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_16 = -1.6562e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_16 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 017, W = 3.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__tvoff_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_17 = 20928.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_17 = -0.0075233
+ sky130_fd_pr__nfet_01v8__pdits_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_17 = 1.513
+ sky130_fd_pr__nfet_01v8__u0_diff_17 = -0.0032502
+ sky130_fd_pr__nfet_01v8__ags_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_17 = 0.001048
+ sky130_fd_pr__nfet_01v8__ua_diff_17 = 1.4247e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_17 = -7.6987e-20
*
* sky130_fd_pr__nfet_01v8, Bin 018, W = 3.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__ub_diff_18 = -1.4311e-20
+ sky130_fd_pr__nfet_01v8__tvoff_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_18 = 9237.1
+ sky130_fd_pr__nfet_01v8__vth0_diff_18 = -0.0029364
+ sky130_fd_pr__nfet_01v8__pdits_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_18 = 1.054
+ sky130_fd_pr__nfet_01v8__u0_diff_18 = -0.0013803
+ sky130_fd_pr__nfet_01v8__ags_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_18 = 0.0023213
+ sky130_fd_pr__nfet_01v8__ua_diff_18 = 3.3268e-12
+ sky130_fd_pr__nfet_01v8__eta0_diff_18 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 019, W = 5.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__eta0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__ua_diff_19 = 2.9314e-12
+ sky130_fd_pr__nfet_01v8__ub_diff_19 = 5.2293e-21
+ sky130_fd_pr__nfet_01v8__tvoff_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_19 = 0.0073134
+ sky130_fd_pr__nfet_01v8__rdsw_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_19 = 0.0012907
+ sky130_fd_pr__nfet_01v8__pdits_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_19 = 0.97435
+ sky130_fd_pr__nfet_01v8__u0_diff_19 = -0.00089361
+ sky130_fd_pr__nfet_01v8__ags_diff_19 = -0.074135
+ sky130_fd_pr__nfet_01v8__keta_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_19 = 0.0053264
*
* sky130_fd_pr__nfet_01v8, Bin 020, W = 5.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__ua_diff_20 = 1.4457e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_20 = -4.6997e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_20 = 0.10627
+ sky130_fd_pr__nfet_01v8__rdsw_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_20 = -0.01318
+ sky130_fd_pr__nfet_01v8__pdits_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_20 = 0.98486
+ sky130_fd_pr__nfet_01v8__u0_diff_20 = -0.0051351
+ sky130_fd_pr__nfet_01v8__ags_diff_20 = -0.05882
+ sky130_fd_pr__nfet_01v8__keta_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_20 = 0.0041307
*
* sky130_fd_pr__nfet_01v8, Bin 021, W = 5.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__ags_diff_21 = -0.085086
+ sky130_fd_pr__nfet_01v8__keta_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_21 = 0.0037858
+ sky130_fd_pr__nfet_01v8__ua_diff_21 = 9.5141e-12
+ sky130_fd_pr__nfet_01v8__eta0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_21 = -3.6045e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_21 = 0.11433
+ sky130_fd_pr__nfet_01v8__rdsw_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_21 = -0.012328
+ sky130_fd_pr__nfet_01v8__pdits_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_21 = 0.92412
+ sky130_fd_pr__nfet_01v8__u0_diff_21 = -0.0036871
*
* sky130_fd_pr__nfet_01v8, Bin 022, W = 5.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__pclm_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_22 = 0.7515
+ sky130_fd_pr__nfet_01v8__u0_diff_22 = -0.0020259
+ sky130_fd_pr__nfet_01v8__ags_diff_22 = -0.024684
+ sky130_fd_pr__nfet_01v8__keta_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_22 = 0.0040638
+ sky130_fd_pr__nfet_01v8__ua_diff_22 = 5.1254e-12
+ sky130_fd_pr__nfet_01v8__eta0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_22 = -1.5425e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_22 = 0.048637
+ sky130_fd_pr__nfet_01v8__rdsw_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_22 = -0.0032552
+ sky130_fd_pr__nfet_01v8__pdits_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_22 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 023, W = 5.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__pditsd_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_23 = 1.2581
+ sky130_fd_pr__nfet_01v8__u0_diff_23 = 0.0017899
+ sky130_fd_pr__nfet_01v8__ags_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_23 = -0.016888
+ sky130_fd_pr__nfet_01v8__ua_diff_23 = -1.1948e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_23 = 1.7359e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_23 = 20779.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_23 = 0.040098
+ sky130_fd_pr__nfet_01v8__pdits_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_23 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 024, W = 5.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__pdits_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_24 = 1.6876
+ sky130_fd_pr__nfet_01v8__u0_diff_24 = -0.0059564
+ sky130_fd_pr__nfet_01v8__ags_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_24 = -0.0064709
+ sky130_fd_pr__nfet_01v8__ua_diff_24 = 4.34e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_24 = -4.6585e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_24 = 12451.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_24 = 0.0060337
+ sky130_fd_pr__nfet_01v8__b0_diff_24 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 025, W = 5.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__b0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_25 = 1.409
+ sky130_fd_pr__nfet_01v8__u0_diff_25 = -0.0027324
+ sky130_fd_pr__nfet_01v8__ags_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_25 = -0.00059331
+ sky130_fd_pr__nfet_01v8__ua_diff_25 = 1.4768e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_25 = 1.8263e-20
+ sky130_fd_pr__nfet_01v8__tvoff_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_25 = 14753.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_25 = 0.0055231
*
* sky130_fd_pr__nfet_01v8, Bin 026, W = 5.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__kt1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_26 = 777.46
+ sky130_fd_pr__nfet_01v8__vth0_diff_26 = 0.0032119
+ sky130_fd_pr__nfet_01v8__b0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_26 = 1.1891
+ sky130_fd_pr__nfet_01v8__u0_diff_26 = -0.00026917
+ sky130_fd_pr__nfet_01v8__ags_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_26 = 0.0022612
+ sky130_fd_pr__nfet_01v8__ua_diff_26 = -3.5035e-13
+ sky130_fd_pr__nfet_01v8__eta0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_26 = 6.1214e-21
+ sky130_fd_pr__nfet_01v8__tvoff_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_26 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 027, W = 7.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__a0_diff_27 = 0.12825
+ sky130_fd_pr__nfet_01v8__rdsw_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_27 = -0.014597
+ sky130_fd_pr__nfet_01v8__b0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_27 = 1.0023
+ sky130_fd_pr__nfet_01v8__u0_diff_27 = -0.002
+ sky130_fd_pr__nfet_01v8__ags_diff_27 = -0.11111
+ sky130_fd_pr__nfet_01v8__keta_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_27 = 0.003022
+ sky130_fd_pr__nfet_01v8__ua_diff_27 = 6.9614e-12
+ sky130_fd_pr__nfet_01v8__eta0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_27 = -8.734e-20
+ sky130_fd_pr__nfet_01v8__tvoff_diff_27 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 028, W = 7.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__tvoff_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_28 = 0.12443
+ sky130_fd_pr__nfet_01v8__rdsw_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_28 = -0.0087303
+ sky130_fd_pr__nfet_01v8__pdits_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_28 = 0.98082
+ sky130_fd_pr__nfet_01v8__u0_diff_28 = -0.0025919
+ sky130_fd_pr__nfet_01v8__ags_diff_28 = -0.086809
+ sky130_fd_pr__nfet_01v8__keta_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_28 = 0.004451
+ sky130_fd_pr__nfet_01v8__ua_diff_28 = 7.1735e-12
+ sky130_fd_pr__nfet_01v8__eta0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_28 = -1.9301e-19
*
* sky130_fd_pr__nfet_01v8, Bin 029, W = 7.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__ub_diff_29 = -1.6863e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_29 = 0.027455
+ sky130_fd_pr__nfet_01v8__rdsw_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_29 = -0.010883
+ sky130_fd_pr__nfet_01v8__pdits_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_29 = 0.90987
+ sky130_fd_pr__nfet_01v8__u0_diff_29 = -0.0023625
+ sky130_fd_pr__nfet_01v8__ags_diff_29 = -0.0070212
+ sky130_fd_pr__nfet_01v8__keta_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_29 = 0.0030976
+ sky130_fd_pr__nfet_01v8__ua_diff_29 = 6.1862e-12
+ sky130_fd_pr__nfet_01v8__eta0_diff_29 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 030, W = 7.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__eta0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_30 = -1.4981e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_30 = 0.06376
+ sky130_fd_pr__nfet_01v8__rdsw_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_30 = -0.0049999
+ sky130_fd_pr__nfet_01v8__pdits_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_30 = 0.88257
+ sky130_fd_pr__nfet_01v8__u0_diff_30 = -0.0019154
+ sky130_fd_pr__nfet_01v8__ags_diff_30 = -0.036504
+ sky130_fd_pr__nfet_01v8__keta_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_30 = 0.0044208
+ sky130_fd_pr__nfet_01v8__ua_diff_30 = 4.8432e-12
*
* sky130_fd_pr__nfet_01v8, Bin 031, W = 7.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__ua_diff_31 = 7.4833e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_31 = 2.652e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_31 = 17673.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_31 = 0.038467
+ sky130_fd_pr__nfet_01v8__pdits_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_31 = -0.73916
+ sky130_fd_pr__nfet_01v8__u0_diff_31 = 0.0037678
+ sky130_fd_pr__nfet_01v8__ags_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_31 = -0.022293
*
* sky130_fd_pr__nfet_01v8, Bin 032, W = 7.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__ags_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_32 = -0.008167
+ sky130_fd_pr__nfet_01v8__ua_diff_32 = 3.5581e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_32 = -3.1684e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_32 = 14059.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_32 = 0.0026594
+ sky130_fd_pr__nfet_01v8__pdits_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_32 = 1.6049
+ sky130_fd_pr__nfet_01v8__u0_diff_32 = -0.0047061
*
* sky130_fd_pr__nfet_01v8, Bin 033, W = 7.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__pclm_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_33 = 1.3243
+ sky130_fd_pr__nfet_01v8__u0_diff_33 = -0.0029225
+ sky130_fd_pr__nfet_01v8__ags_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_33 = -0.00069916
+ sky130_fd_pr__nfet_01v8__ua_diff_33 = 1.7019e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_33 = -1.0021e-20
+ sky130_fd_pr__nfet_01v8__tvoff_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_33 = 16966.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_33 = 0.00050461
+ sky130_fd_pr__nfet_01v8__pdits_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_33 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 034, W = 7.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8__pditsd_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_34 = 1.1492
+ sky130_fd_pr__nfet_01v8__u0_diff_34 = -0.00026741
+ sky130_fd_pr__nfet_01v8__ags_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_34 = 0.0014281
+ sky130_fd_pr__nfet_01v8__ua_diff_34 = -2.9115e-13
+ sky130_fd_pr__nfet_01v8__eta0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_34 = -1.225e-20
+ sky130_fd_pr__nfet_01v8__tvoff_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_34 = 1851.3
+ sky130_fd_pr__nfet_01v8__kt1_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_34 = 0.00010691
+ sky130_fd_pr__nfet_01v8__pdits_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_34 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 035, W = 0.42u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__pdits_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_35 = 1.6547e-8
+ sky130_fd_pr__nfet_01v8__pditsd_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_35 = 1.4052
+ sky130_fd_pr__nfet_01v8__u0_diff_35 = -0.009592
+ sky130_fd_pr__nfet_01v8__ags_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_35 = 0.00133
+ sky130_fd_pr__nfet_01v8__ua_diff_35 = 2.5805e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_35 = -4.365e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_35 = 0.0091492
+ sky130_fd_pr__nfet_01v8__b0_diff_35 = -2.2934e-7
*
* sky130_fd_pr__nfet_01v8, Bin 036, W = 0.42u, L = 20.0u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__b0_diff_36 = 1.7766e-11
+ sky130_fd_pr__nfet_01v8__pdits_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_36 = 1.0478e-8
+ sky130_fd_pr__nfet_01v8__pditsd_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_36 = 2.0416
+ sky130_fd_pr__nfet_01v8__u0_diff_36 = -0.0067261
+ sky130_fd_pr__nfet_01v8__ags_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_36 = 0.0087245
+ sky130_fd_pr__nfet_01v8__ua_diff_36 = 1.5099e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_36 = -4.0381e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_36 = -0.015174
*
* sky130_fd_pr__nfet_01v8, Bin 037, W = 0.42u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__kt1_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_37 = -0.025738
+ sky130_fd_pr__nfet_01v8__b0_diff_37 = -2.5484e-8
+ sky130_fd_pr__nfet_01v8__pdits_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_37 = 2.2209e-8
+ sky130_fd_pr__nfet_01v8__pditsd_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_37 = 1.2926
+ sky130_fd_pr__nfet_01v8__u0_diff_37 = -0.01
+ sky130_fd_pr__nfet_01v8__ags_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_37 = 0.0040008
+ sky130_fd_pr__nfet_01v8__ua_diff_37 = 5.0068e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_37 = -5.9906e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_37 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 038, W = 0.42u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__a0_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_38 = -0.019101
+ sky130_fd_pr__nfet_01v8__b0_diff_38 = -3.2922e-8
+ sky130_fd_pr__nfet_01v8__pdits_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_38 = 9.7406e-9
+ sky130_fd_pr__nfet_01v8__pditsd_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_38 = 1.2083
+ sky130_fd_pr__nfet_01v8__u0_diff_38 = -0.0067325
+ sky130_fd_pr__nfet_01v8__ags_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_38 = 0.0080533
+ sky130_fd_pr__nfet_01v8__ua_diff_38 = 1.7212e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_38 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_38 = -3.8713e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_38 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 039, W = 0.42u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__tvoff_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_39 = -0.0064501
+ sky130_fd_pr__nfet_01v8__pdits_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_39 = 1.7542e-8
+ sky130_fd_pr__nfet_01v8__b1_diff_39 = 8.3616e-9
+ sky130_fd_pr__nfet_01v8__pditsd_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_39 = 1.651
+ sky130_fd_pr__nfet_01v8__u0_diff_39 = -0.0067958
+ sky130_fd_pr__nfet_01v8__ags_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_39 = 0.0015739
+ sky130_fd_pr__nfet_01v8__ua_diff_39 = 1.5825e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_39 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_39 = -4.5424e-19
*
* sky130_fd_pr__nfet_01v8, Bin 040, W = 0.42u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__tvoff_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_40 = 65211.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_40 = 0.06351
+ sky130_fd_pr__nfet_01v8__pdits_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_40 = 0.58732
+ sky130_fd_pr__nfet_01v8__u0_diff_40 = -0.0040023
+ sky130_fd_pr__nfet_01v8__ags_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_40 = -0.015063
+ sky130_fd_pr__nfet_01v8__ua_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__eta0_diff_40 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_40 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 041, W = 0.42u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__eta0_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_41 = -7.3036e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_41 = 31134.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_41 = 0.0079464
+ sky130_fd_pr__nfet_01v8__pdits_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_41 = -0.40516
+ sky130_fd_pr__nfet_01v8__u0_diff_41 = -0.01086
+ sky130_fd_pr__nfet_01v8__ags_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_41 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_41 = -0.010225
+ sky130_fd_pr__nfet_01v8__ua_diff_41 = 4.5834e-11
*
* sky130_fd_pr__nfet_01v8, Bin 042, W = 0.42u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__ua_diff_42 = 5.2591e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_42 = -4.2543e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_42 = 100000.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_42 = 0.019407
+ sky130_fd_pr__nfet_01v8__pdits_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_42 = -0.040061
+ sky130_fd_pr__nfet_01v8__b1_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_42 = -0.01641
+ sky130_fd_pr__nfet_01v8__u0_diff_42 = -0.0080919
+ sky130_fd_pr__nfet_01v8__ags_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_42 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_42 = 0.0064036
*
* sky130_fd_pr__nfet_01v8, Bin 043, W = 0.55u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__ags_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_43 = 0.003968
+ sky130_fd_pr__nfet_01v8__ua_diff_43 = 1.7661e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_43 = -2.786e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_43 = 0.016392
+ sky130_fd_pr__nfet_01v8__pdits_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_43 = 8.0476e-8
+ sky130_fd_pr__nfet_01v8__voff_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_43 = 1.1223e-8
+ sky130_fd_pr__nfet_01v8__pditsd_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_43 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_43 = 1.1484
+ sky130_fd_pr__nfet_01v8__u0_diff_43 = -0.0064337
*
* sky130_fd_pr__nfet_01v8, Bin 044, W = 0.55u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__pclm_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_44 = 1.4963
+ sky130_fd_pr__nfet_01v8__u0_diff_44 = -0.01
+ sky130_fd_pr__nfet_01v8__ags_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_44 = 0.007003
+ sky130_fd_pr__nfet_01v8__ua_diff_44 = 1.4279e-10
+ sky130_fd_pr__nfet_01v8__eta0_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_44 = -9.0211e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_44 = -0.013358
+ sky130_fd_pr__nfet_01v8__pdits_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_44 = 2.0197e-8
+ sky130_fd_pr__nfet_01v8__voff_diff_44 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_44 = 2.1661e-8
+ sky130_fd_pr__nfet_01v8__pditsd_diff_44 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 045, W = 0.55u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__pditsd_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_45 = 0.95211
+ sky130_fd_pr__nfet_01v8__u0_diff_45 = -0.0067575
+ sky130_fd_pr__nfet_01v8__ags_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_45 = 0.0018992
+ sky130_fd_pr__nfet_01v8__ua_diff_45 = 1.8192e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_45 = -4.3254e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_45 = -0.0029178
+ sky130_fd_pr__nfet_01v8__pdits_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_45 = -6.9109e-9
+ sky130_fd_pr__nfet_01v8__voff_diff_45 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_45 = 7.9176e-9
*
* sky130_fd_pr__nfet_01v8, Bin 046, W = 0.55u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__pdits_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_46 = 8.4769e-9
+ sky130_fd_pr__nfet_01v8__pditsd_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_46 = 1.4216
+ sky130_fd_pr__nfet_01v8__u0_diff_46 = -0.0050966
+ sky130_fd_pr__nfet_01v8__ags_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_46 = 0.0054045
+ sky130_fd_pr__nfet_01v8__ua_diff_46 = 1.3113e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_46 = -2.2805e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_46 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_46 = -0.0028103
+ sky130_fd_pr__nfet_01v8__b0_diff_46 = 2.6687e-9
*
* sky130_fd_pr__nfet_01v8, Bin 047, W = 0.55u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__b0_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_47 = -0.014371
+ sky130_fd_pr__nfet_01v8__b1_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_47 = -0.4183
+ sky130_fd_pr__nfet_01v8__u0_diff_47 = -0.0021722
+ sky130_fd_pr__nfet_01v8__ags_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_47 = -0.016152
+ sky130_fd_pr__nfet_01v8__ua_diff_47 = 1.5346e-10
+ sky130_fd_pr__nfet_01v8__eta0_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_47 = 1.6496e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_47 = 100000.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_47 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_47 = 0.063549
*
* sky130_fd_pr__nfet_01v8, Bin 048, W = 0.55u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__kt1_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_48 = 39250.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_48 = 0.0073028
+ sky130_fd_pr__nfet_01v8__b0_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_48 = 1.7187
+ sky130_fd_pr__nfet_01v8__u0_diff_48 = -0.0053846
+ sky130_fd_pr__nfet_01v8__ags_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_48 = 0.0027652
+ sky130_fd_pr__nfet_01v8__ua_diff_48 = 1.1686e-11
+ sky130_fd_pr__nfet_01v8__eta0_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_48 = -3.1734e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_48 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_48 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 049, W = 0.64u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__a0_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_49 = 37983.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_49 = 0.079991
+ sky130_fd_pr__nfet_01v8__b0_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_49 = 0.22483
+ sky130_fd_pr__nfet_01v8__u0_diff_49 = -0.0038167
+ sky130_fd_pr__nfet_01v8__ags_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_49 = -0.015958
+ sky130_fd_pr__nfet_01v8__ua_diff_49 = 1.3513e-10
+ sky130_fd_pr__nfet_01v8__eta0_diff_49 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_49 = -5.5497e-19
+ sky130_fd_pr__nfet_01v8__tvoff_diff_49 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 050, W = 0.84u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__tvoff_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_50 = 56151.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_50 = 0.048934
+ sky130_fd_pr__nfet_01v8__pdits_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__nfactor_diff_50 = 0.22447
+ sky130_fd_pr__nfet_01v8__u0_diff_50 = -0.0023891
+ sky130_fd_pr__nfet_01v8__ags_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__keta_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_50 = -0.017649
+ sky130_fd_pr__nfet_01v8__ua_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__eta0_diff_50 = 0.0
+ sky130_fd_pr__nfet_01v8__ub_diff_50 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 051, W = 0.74u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__tvoff_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_51 = 44079.09414086
+ sky130_fd_pr__nfet_01v8__kt1_diff_51 = -4.96639e-5
+ sky130_fd_pr__nfet_01v8__vth0_diff_51 = 0.06735546
+ sky130_fd_pr__nfet_01v8__pdits_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_51 = -0.00027261
+ sky130_fd_pr__nfet_01v8__u0_diff_51 = -0.00019859
+ sky130_fd_pr__nfet_01v8__nfactor_diff_51 = -0.15794521
+ sky130_fd_pr__nfet_01v8__keta_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_51 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_51 = -0.01908401
+ sky130_fd_pr__nfet_01v8__ua_diff_51 = 4.61938e-11
+ sky130_fd_pr__nfet_01v8__ub_diff_51 = -1.76062e-19
+ sky130_fd_pr__nfet_01v8__eta0_diff_51 = -6.59195e-17
*
* sky130_fd_pr__nfet_01v8, Bin 052, W = 0.36u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__ub_diff_52 = -1.32884e-18
+ sky130_fd_pr__nfet_01v8__eta0_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__tvoff_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_52 = 31459.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_52 = 0.14691
+ sky130_fd_pr__nfet_01v8__pdits_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_52 = 0.0112789
+ sky130_fd_pr__nfet_01v8__pditsd_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_52 = -0.00090237
+ sky130_fd_pr__nfet_01v8__u0_diff_52 = -0.017871
+ sky130_fd_pr__nfet_01v8__nfactor_diff_52 = 0.55976134
+ sky130_fd_pr__nfet_01v8__keta_diff_52 = -0.00301097
+ sky130_fd_pr__nfet_01v8__ags_diff_52 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_52 = 0.0084041
+ sky130_fd_pr__nfet_01v8__ua_diff_52 = -9.72898e-11
*
* sky130_fd_pr__nfet_01v8, Bin 053, W = 0.39u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__ua_diff_53 = -4.01828e-11
+ sky130_fd_pr__nfet_01v8__ub_diff_53 = -9.60681e-19
+ sky130_fd_pr__nfet_01v8__eta0_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__tvoff_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_53 = 37070.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_53 = 0.13857
+ sky130_fd_pr__nfet_01v8__pdits_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_53 = 0.00507783
+ sky130_fd_pr__nfet_01v8__pditsd_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_53 = -0.00031247
+ sky130_fd_pr__nfet_01v8__u0_diff_53 = -0.012893
+ sky130_fd_pr__nfet_01v8__nfactor_diff_53 = 0.17556582
+ sky130_fd_pr__nfet_01v8__keta_diff_53 = -0.00104263
+ sky130_fd_pr__nfet_01v8__ags_diff_53 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_53 = 0.00316
*
* sky130_fd_pr__nfet_01v8, Bin 054, W = 0.52u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__keta_diff_54 = 0.00033095
+ sky130_fd_pr__nfet_01v8__ags_diff_54 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_54 = -0.015566
+ sky130_fd_pr__nfet_01v8__ua_diff_54 = 1.14081e-10
+ sky130_fd_pr__nfet_01v8__ub_diff_54 = 7.22805e-20
+ sky130_fd_pr__nfet_01v8__eta0_diff_54 = 3.51265e-6
+ sky130_fd_pr__nfet_01v8__tvoff_diff_54 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_54 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_54 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_54 = 129550.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_54 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_54 = 0.10173
+ sky130_fd_pr__nfet_01v8__pdits_diff_54 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_54 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_54 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_54 = -0.01182365
+ sky130_fd_pr__nfet_01v8__pditsd_diff_54 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_54 = 9.91854e-5
+ sky130_fd_pr__nfet_01v8__u0_diff_54 = -0.0021466
+ sky130_fd_pr__nfet_01v8__nfactor_diff_54 = -0.89046554
*
* sky130_fd_pr__nfet_01v8, Bin 055, W = 0.54u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__pclm_diff_55 = 3.63878e-5
+ sky130_fd_pr__nfet_01v8__u0_diff_55 = -0.00011811
+ sky130_fd_pr__nfet_01v8__nfactor_diff_55 = -1.00161089
+ sky130_fd_pr__nfet_01v8__keta_diff_55 = 0.00012142
+ sky130_fd_pr__nfet_01v8__ags_diff_55 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_55 = -0.016319
+ sky130_fd_pr__nfet_01v8__ua_diff_55 = 1.29803e-10
+ sky130_fd_pr__nfet_01v8__ub_diff_55 = 1.80964e-19
+ sky130_fd_pr__nfet_01v8__eta0_diff_55 = 1.28866e-6
+ sky130_fd_pr__nfet_01v8__tvoff_diff_55 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_55 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_55 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_55 = 114670.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_55 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_55 = 0.098686
+ sky130_fd_pr__nfet_01v8__pdits_diff_55 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_55 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_55 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_55 = -0.01355952
+ sky130_fd_pr__nfet_01v8__pditsd_diff_55 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 056, W = 0.58u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__pditsd_diff_56 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_56 = 6.70187e-5
+ sky130_fd_pr__nfet_01v8__u0_diff_56 = -0.0020688
+ sky130_fd_pr__nfet_01v8__nfactor_diff_56 = -0.75172882
+ sky130_fd_pr__nfet_01v8__keta_diff_56 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_56 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_56 = -0.016241
+ sky130_fd_pr__nfet_01v8__ua_diff_56 = 1.32078e-10
+ sky130_fd_pr__nfet_01v8__ub_diff_56 = -1.42771e-20
+ sky130_fd_pr__nfet_01v8__eta0_diff_56 = -2.37352e-6
+ sky130_fd_pr__nfet_01v8__tvoff_diff_56 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_56 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_56 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_56 = 117840.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_56 = 3.41931e-5
+ sky130_fd_pr__nfet_01v8__vth0_diff_56 = 0.096363
+ sky130_fd_pr__nfet_01v8__pdits_diff_56 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_56 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_56 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_56 = -0.00899558
*
* sky130_fd_pr__nfet_01v8, Bin 057, W = 0.6u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__pdits_diff_57 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_57 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_57 = -0.00576244
+ sky130_fd_pr__nfet_01v8__pditsd_diff_57 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_57 = 6.89796e-5
+ sky130_fd_pr__nfet_01v8__u0_diff_57 = -0.0033469
+ sky130_fd_pr__nfet_01v8__nfactor_diff_57 = -0.56979137
+ sky130_fd_pr__nfet_01v8__keta_diff_57 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_57 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_57 = -0.01636
+ sky130_fd_pr__nfet_01v8__ua_diff_57 = 1.2904e-10
+ sky130_fd_pr__nfet_01v8__ub_diff_57 = -1.61883e-19
+ sky130_fd_pr__nfet_01v8__eta0_diff_57 = -2.44296e-6
+ sky130_fd_pr__nfet_01v8__tvoff_diff_57 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_57 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_57 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_57 = 131300.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_57 = 3.51936e-5
+ sky130_fd_pr__nfet_01v8__vth0_diff_57 = 0.093492
+ sky130_fd_pr__nfet_01v8__b0_diff_57 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 058, W = 0.61u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__b0_diff_58 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_58 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_58 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_58 = -0.00423892
+ sky130_fd_pr__nfet_01v8__pditsd_diff_58 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_58 = 5.98153e-5
+ sky130_fd_pr__nfet_01v8__u0_diff_58 = -0.0035976
+ sky130_fd_pr__nfet_01v8__nfactor_diff_58 = -0.48397308
+ sky130_fd_pr__nfet_01v8__keta_diff_58 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_58 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_58 = -0.016314
+ sky130_fd_pr__nfet_01v8__ua_diff_58 = 1.27611e-10
+ sky130_fd_pr__nfet_01v8__ub_diff_58 = -2.3131e-19
+ sky130_fd_pr__nfet_01v8__eta0_diff_58 = -2.11841e-6
+ sky130_fd_pr__nfet_01v8__tvoff_diff_58 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_58 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_58 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_58 = 117490.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_58 = 3.05179e-5
+ sky130_fd_pr__nfet_01v8__vth0_diff_58 = 0.092388
*
* sky130_fd_pr__nfet_01v8, Bin 059, W = 0.65u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__kt1_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_59 = 68805.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_59 = 0.090402
+ sky130_fd_pr__nfet_01v8__b0_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__pdits_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_59 = -6.90229e-5
+ sky130_fd_pr__nfet_01v8__u0_diff_59 = -0.0052071
+ sky130_fd_pr__nfet_01v8__nfactor_diff_59 = -0.23492281
+ sky130_fd_pr__nfet_01v8__keta_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_59 = -0.016096
+ sky130_fd_pr__nfet_01v8__ua_diff_59 = 1.14656e-10
+ sky130_fd_pr__nfet_01v8__ub_diff_59 = -3.9518e-19
+ sky130_fd_pr__nfet_01v8__eta0_diff_59 = 2.82807e-17
+ sky130_fd_pr__nfet_01v8__tvoff_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_59 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_59 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 060, W = 0.65u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__vsat_diff_60 = 58947.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_60 = 0.06508
+ sky130_fd_pr__nfet_01v8__pdits_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_60 = -6.90233e-5
+ sky130_fd_pr__nfet_01v8__u0_diff_60 = -0.0032164
+ sky130_fd_pr__nfet_01v8__nfactor_diff_60 = -0.23492281
+ sky130_fd_pr__nfet_01v8__keta_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_60 = -0.0081138
+ sky130_fd_pr__nfet_01v8__ua_diff_60 = 1.14656e-10
+ sky130_fd_pr__nfet_01v8__ub_diff_60 = -3.9518e-19
+ sky130_fd_pr__nfet_01v8__eta0_diff_60 = 2.41337e-11
+ sky130_fd_pr__nfet_01v8__tvoff_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_60 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_60 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 061, W = 0.65u, L = 0.25u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8__tvoff_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_61 = 55439.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_61 = 0.027531
+ sky130_fd_pr__nfet_01v8__pdits_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__b1_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__voff_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__u0_diff_61 = -0.0063455
+ sky130_fd_pr__nfet_01v8__nfactor_diff_61 = -0.37468
+ sky130_fd_pr__nfet_01v8__keta_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_61 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_61 = -0.0044406
+ sky130_fd_pr__nfet_01v8__ua_diff_61 = 6.2172e-11
+ sky130_fd_pr__nfet_01v8__ub_diff_61 = -6.17181e-19
+ sky130_fd_pr__nfet_01v8__eta0_diff_61 = 0.0
*
* sky130_fd_pr__nfet_01v8, Bin 062, W = 0.65u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8__tvoff_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__rdsw_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__a0_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__vsat_diff_62 = 99416.0
+ sky130_fd_pr__nfet_01v8__kt1_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__vth0_diff_62 = 0.02186
+ sky130_fd_pr__nfet_01v8__pdits_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__b0_diff_62 = -4.12989e-17
+ sky130_fd_pr__nfet_01v8__b1_diff_62 = 6.53778e-18
+ sky130_fd_pr__nfet_01v8__voff_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__pditsd_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__pclm_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__u0_diff_62 = -0.0035194
+ sky130_fd_pr__nfet_01v8__nfactor_diff_62 = 0.0618
+ sky130_fd_pr__nfet_01v8__keta_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__ags_diff_62 = 0.0
+ sky130_fd_pr__nfet_01v8__k2_diff_62 = 0.0019275
+ sky130_fd_pr__nfet_01v8__ua_diff_62 = 7.7528e-12
+ sky130_fd_pr__nfet_01v8__ub_diff_62 = -3.1358e-19
+ sky130_fd_pr__nfet_01v8__eta0_diff_62 = 0.0
*.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_01v8.pm3.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_01v8__ss.pm3.spice"
