* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 11
.param
+ sky130_fd_pr__nfet_05v0_nvt__toxe_mult = 0.9635
+ sky130_fd_pr__nfet_05v0_nvt__rshn_mult = 1.0
+ sky130_fd_pr__nfet_05v0_nvt__overlap_mult = 5.1025e-1
+ sky130_fd_pr__nfet_05v0_nvt__ajunction_mult = 6.8772e-1
+ sky130_fd_pr__nfet_05v0_nvt__pjunction_mult = 9.0190e-1
+ sky130_fd_pr__nfet_05v0_nvt__lint_diff = 1.21275e-8
+ sky130_fd_pr__nfet_05v0_nvt__wint_diff = -2.252e-8
+ sky130_fd_pr__nfet_05v0_nvt__dlc_diff = 1.6112e-8
+ sky130_fd_pr__nfet_05v0_nvt__dwc_diff = -2.252e-8
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 000, W = 10.0u, L = 2.0u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_0 = 0.056665
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_0 = -0.052927
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_0 = -0.00059672
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_0 = -0.0090633
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_0 = -3.141e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_0 = -0.030851
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_0 = -0.005637
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_0 = -1.5907e-18
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 001, W = 10.0u, L = 4.0u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_1 = -1.357e-18
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_1 = -0.019967
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_1 = -0.032965
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_1 = -0.0051327
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_1 = -0.0077525
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_1 = -2.636e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_1 = -0.018137
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_1 = -0.0051202
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 002, W = 10.0u, L = 0.9u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_2 = -1.8782e-18
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_2 = 0.066292
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_2 = 0.00087158
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_2 = -0.0096682
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_2 = -4.2384e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_2 = -6160.2
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_2 = -0.03046
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_2 = 0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 003, W = 1.0u, L = 25.0u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_3 = -2.0373e-11
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_3 = -0.0020789
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_3 = -1.0928e-18
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_3 = 0.015653
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_3 = 0.0012297
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_3 = -0.0052343
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_3 = -0.0065532
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_3 = -0.024011
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 004, W = 1.0u, L = 2.0u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_4 = -0.0083037
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_4 = -0.020154
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_4 = -2.6021e-11
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_4 = -0.038115
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_4 = -1.4421e-18
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_4 = -0.05753
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_4 = -0.17718
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_4 = -0.0022264
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 005, W = 1.0u, L = 4.0u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_5 = -0.00093844
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_5 = -0.007664
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_5 = -0.017363
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_5 = -2.4895e-11
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_5 = -0.0093971
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_5 = -1.3242e-18
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_5 = -0.0035696
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_5 = -0.044469
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_5 = 0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 006, W = 1.0u, L = 8.0u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_6 = -0.047321
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_6 = -0.0028201
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_6 = -0.0068477
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_6 = -0.023509
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_6 = -2.2313e-11
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_6 = -0.009358
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_6 = -1.1832e-18
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_6 = -0.022424
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 007, W = 1.0u, L = 0.9u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_7 = 0.043963
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_7 = -3.5325e-6
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_7 = -0.010425
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_7 = -0.038579
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_7 = -3.6456e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_7 = -6428.9
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_7 = -1.7165e-18
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_7 = 0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 008, W = 0.42u, L = 1.0u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_8 = 0.017354
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_8 = 1.5203e-7
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_8 = -0.0095342
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_8 = -0.0085304
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_8 = -0.055166
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_8 = -3.4036e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_8 = -4.5502e-9
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_8 = -1.6434e-18
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_8 = 0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 009, W = 0.42u, L = 0.9u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_9 = -0.13265
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_9 = -0.0070168
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_9 = -0.0087887
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_9 = -0.042098
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_9 = -2.2834e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_9 = -8459.3
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_9 = -1.3613e-18
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 010, W = 0.7u, L = 0.9u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_10 = -7916.1
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_10 = -0.035797
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_10 = 0.028686
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_10 = -0.010001
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_10 = 0.00041829
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_10 = -3.5554e-11
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_10 = -1.6633e-18
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_10 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_05v0_nvt.pm3.spice"
