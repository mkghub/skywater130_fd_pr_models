* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 18
.param
+ sky130_fd_pr__rf_pfet_01v8_b__toxe_mult = 0.948
+ sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult = 0.8
+ sky130_fd_pr__rf_pfet_01v8_b__overlap_mult = 0.95436
+ sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult = 0.90161
+ sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult = 0.90587
+ sky130_fd_pr__rf_pfet_01v8_b__lint_diff = 1.7325e-8
+ sky130_fd_pr__rf_pfet_01v8_b__wint_diff = -3.2175e-8
+ sky130_fd_pr__rf_pfet_01v8_b__rshg_diff = -7.0
+ sky130_fd_pr__rf_pfet_01v8_b__xgw_diff = -6.425e-8
+ sky130_fd_pr__rf_pfet_01v8_b__dlc_diff = 1.7325e-8
+ sky130_fd_pr__rf_pfet_01v8_b__dwc_diff = 0.0
+ sky130_fd_pr__rf_pfet_01v8__aw_cap_mult = 0.85
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult = 0.77
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult = 0.77
+ sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2 = 0.85
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2 = 0.80
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2 = 0.80
+ sky130_fd_pr__rf_pfet_01v8__aw_rd_mult = 1.0
+ sky130_fd_pr__rf_pfet_01v8__aw_rs_mult = 1.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_0 = 0.0036576
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_0 = -0.00034614
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_0 = -0.09351
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_0 = -19636.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_0 = -0.39184
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_0 = 0.53599
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_0 = -0.0076131
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_0 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_1 = -0.0076806
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_1 = -0.00019683
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_1 = -0.08358
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_1 = -15546.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_1 = -0.55481
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_1 = 0.94783
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_1 = -0.10922
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_1 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_2 = -0.15
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_2 = -0.033345
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_2 = -3.0791e-5
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_2 = 0.00085561
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_2 = -6434.1
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_2 = -0.73688
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_2 = 5.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_2 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_3 = 0.039133
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_3 = -0.0012925
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_3 = -0.00028011
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_3 = -0.11455
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_3 = -18686.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_3 = -0.31125
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_3 = 0.13079
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_3 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_4 = -0.58068
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_4 = 0.48528
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_4 = -0.051759
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_4 = 0.00024736
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_4 = -0.00041476
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_4 = -0.075262
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_4 = -11333.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_4 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_5 = -0.7435
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_5 = 5.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_5 = -0.15
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_5 = -0.016582
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_5 = -0.00016695
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_5 = -0.0082165
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_5 = -1107.2
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_5 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_6 = -0.37364
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_6 = -0.0015912
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_6 = 0.04821
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_6 = -0.0014721
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_6 = -0.00053506
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_6 = -0.12391
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_6 = -16484.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_7 = -0.00025473
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_7 = -17993.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_7 = -0.49017
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_7 = 0.77211
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_7 = -0.070464
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_7 = 0.00033491
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_7 = -0.084215
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_8 = -0.057631
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_8 = -0.00020922
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_8 = -5719.7
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_8 = -0.6769
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_8 = 4.6157
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_8 = -0.15
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_8 = -0.019564
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_0 = 0.0065905
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_0 = -0.38688
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_0 = -0.19049
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_0 = 0.050397
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_0 = -0.00050702
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_0 = -0.078819
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_0 = -20196.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_1 = -12293.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_1 = -0.0063812
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_1 = -0.43628
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_1 = 0.60205
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_1 = -0.09979
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_1 = -0.00027314
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_1 = -0.068972
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_2 = -7.2735e-5
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_2 = -0.041687
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_2 = 272.66
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_2 = -0.034415
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_2 = -0.65512
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_2 = 5.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_2 = -0.15
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_2 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_3 = 0.055428
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_3 = -0.0003818
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_3 = -0.10701
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_3 = -16139.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_3 = 0.00078898
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_3 = -0.22318
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_3 = 0.31839
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_3 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_4 = -0.031099
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_4 = -0.00058216
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_4 = -0.060108
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_4 = -11485.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_4 = 0.0039762
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_4 = -0.47494
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_4 = 0.23524
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_5 = -0.15
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_5 = -0.04076
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_5 = -0.00025609
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_5 = -7303.4
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_5 = -0.016473
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_5 = -0.59835
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_5 = 4.4656
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_6 = -0.33154
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_6 = -0.15691
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_6 = 0.089833
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_6 = -0.10181
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_6 = -0.00035343
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_6 = -16543.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_6 = 0.00030278
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_7 = 0.0028314
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_7 = -0.41124
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_7 = 0.44953
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_7 = -0.045335
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_7 = -0.077646
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_7 = -0.000511
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_7 = -15224.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_7 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_8 = -0.018202
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_8 = -0.55037
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_8 = 3.1422
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_8 = -0.15
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_8 = -0.037861
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_8 = -0.00030626
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_8 = 4136.5
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_8 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__rf_pfet_01v8_b.pm3.spice"
