* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
*
* model corner
* , Bin 000, W = 30.0u, L = 1.0u
* ----------------------------
.param
+ sky130_fd_pr__nfet_20v0_nvt__rdrift_mult = 1.3479e+0
+ sky130_fd_pr__nfet_20v0_nvt__hvvsat_mult = 7.9823e-1
+ sky130_fd_pr__nfet_20v0_nvt__vth0_diff = 1.6910e-1
+ sky130_fd_pr__nfet_20v0_nvt__k2_diff = -1.1937e-1
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_20v0_nvt__subcircuit.pm3.spice"
