* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 18
.param
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult = 0.9635
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult = 0.8
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult = 8.8119e-1
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult = 8.7784e-1
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult = 7.8244e-1
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff = 1.21275e-8
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff = -2.252e-8
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff = -7.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff = 7.7131e-9
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff = -4.504e-8
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42 = 0.8875
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42 = 0.755
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42 = 0.755
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult = 0.8875
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult = 0.825
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult = 0.825
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult = 1.0
+ sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult = 1.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_0 = -0.043187
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_0 = 0.0031893
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_0 = -20156.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_0 = -0.0091082
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_1 = -0.00023031
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_1 = -0.039728
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_1 = 0.0032163
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_1 = -16799.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_1 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_2 = -0.0031116
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_2 = -0.032085
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_2 = 0.003301
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_2 = -12923.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_2 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_3 = 0.0056278
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_3 = -0.051298
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_3 = -0.001719
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_3 = -25716.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_3 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_4 = 0.0040629
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_4 = -0.050969
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_4 = -0.001606
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_4 = -16982.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_4 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_5 = 0.0028518
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_5 = -0.021748
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_5 = 0.001153
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_5 = -11783.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_5 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_6 = -0.0053048
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_6 = -0.045076
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_6 = -0.0074793
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_6 = -20834.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_6 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_7 = 0.0027467
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_7 = -0.042761
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_7 = -0.0034925
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_7 = -14000.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_7 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__pclm_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__k2_diff_8 = 0.0026278
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vth0_diff_8 = -0.018088
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__u0_diff_8 = 0.00072051
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__vsat_diff_8 = -10215.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM02__b1_diff_8 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_0 = -0.0093685
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_0 = -0.046477
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_0 = -0.003305
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_0 = -16286.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_0 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_1 = -0.0011171
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_1 = -0.047694
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_1 = -0.00091767
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_1 = -16903.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_1 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_2 = 0.0014264
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_2 = -0.037401
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_2 = 0.00086418
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_2 = -7635.6
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_2 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_3 = 0.004034
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_3 = -0.049369
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_3 = -0.0026239
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_3 = -26112.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_4 = -0.0064811
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_4 = -15470.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_4 = 0.002107
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_4 = -0.046682
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_5 = -0.033495
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_5 = -0.002231
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_5 = -2766.3
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_5 = 0.0013838
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_6 = -0.0022088
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_6 = -0.049429
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_6 = -0.0050469
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_6 = -24301.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_6 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_7 = -0.00079282
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_7 = -0.042712
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_7 = -0.0075496
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_7 = -16463.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_7 = 0.0
*
* sky130_fd_pr__rf_nfet_01v8_lvt_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__pclm_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__k2_diff_8 = 0.00082322
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__u0_diff_8 = -0.0041644
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vsat_diff_8 = -543.48
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__vth0_diff_8 = -0.034543
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_nfet_01v8_lvt_bM04__ua_diff_8 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"
