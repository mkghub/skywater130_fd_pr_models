* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 8
.param
+ sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult = 1.06
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult = 1.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult = 1.292
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult = 1.0777e+0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult = 1.0736e+0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff = -1.7325e-8
+ sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff = 3.2175e-8
+ sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff = -1.7325e-8
+ sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff = 3.2175e-8
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 000, W = 14.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_0 = 8.3700e-3
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_0 = 2.6732e-3
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_0 = 9.4633e+4
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_0 = -5.8555e-2
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_0 = -4.2555e-1
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_0 = 1.9037e-10
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_0 = 1.0572e-18
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_0 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_0 = -1.1583e-3
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 001, W = 15.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_1 = 0.15309
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_1 = 0.015841
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_1 = -0.0066616
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_1 = 22080.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_1 = 0.070909
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_1 = -5.5136e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_1 = 0.51452
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_1 = -3.0377e-18
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_1 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_1 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 002, W = 16.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_2 = 5.4092e-2
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_2 = 1.0843e-2
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_2 = 2.4584e-4
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_2 = -2.9721e-2
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_2 = 3.6720e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_2 = 6.4607e+4
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_2 = 3.7549e-1
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_2 = 1.9733e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_2 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_2 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 003, W = 17.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_3 = 3.3063e-2
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_3 = 9.1109e-3
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_3 = 2.0202e-3
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_3 = -5.2973e-2
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_3 = 7.2069e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_3 = 4.3170e+4
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_3 = 1.2833e-1
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_3 = 7.6394e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_3 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_3 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 004, W = 19.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_4 = 0.022785
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_4 = 0.0088938
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_4 = 0.0020785
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_4 = '-0.06018-0.005'
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_4 = 5.9115e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_4 = 47898.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_4 = -0.1672
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_4 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_4 = 9.8318e-19
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_4 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 005, W = 21.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_5 = 0.16248
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_5 = 0.016552
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_5 = -0.0073777
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_5 = 0.078938
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_5 = -5.267e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_5 = 28612.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_5 = 0.56919
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_5 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_5 = -3.3626e-18
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 006, W = 23.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_6 = -3.936e-18
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_6 = 0.18617
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_6 = 0.016075
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_6 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_6 = -0.0087419
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_6 = 0.11079
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_6 = -4.0545e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_6 = 40444.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_6 = 0.47252
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_6 = 0.0
*
* sky130_fd_pr__esd_pfet_g5v0d10v5, Bin 007, W = 26.5u, L = 0.55u
* -----------------------------------
+ sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_7 = -2.7759e-18
+ sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_7 = 0.14442
+ sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_7 = 0.016523
+ sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_7 = 0.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_7 = -0.006295
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_7 = 0.059613
+ sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_7 = 1.6811e-11
+ sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_7 = 21388.0
+ sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_7 = 0.57083
+ sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_7 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice"
