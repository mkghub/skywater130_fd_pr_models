* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 8
.param
+ sky130_fd_pr__rf_pfet_01v8_b__toxe_mult = 1.052
+ sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult = 1.2
+ sky130_fd_pr__rf_pfet_01v8_b__overlap_mult = 1.1934
+ sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult = 1.0909
+ sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult = 1.096
+ sky130_fd_pr__rf_pfet_01v8_b__lint_diff = -1.7325e-8
+ sky130_fd_pr__rf_pfet_01v8_b__wint_diff = 3.2175e-8
+ sky130_fd_pr__rf_pfet_01v8_b__rshg_diff = 7.0
+ sky130_fd_pr__rf_pfet_01v8_b__dlc_diff = -1.7325e-8
+ sky130_fd_pr__rf_pfet_01v8_b__dwc_diff = 0.0
+ sky130_fd_pr__rf_pfet_01v8_b__xgw_diff = 6.4250e-8
+ sky130_fd_pr__rf_pfet_01v8__aw_cap_mult = 1.15
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult = 1.45
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult = 1.45
+ sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2 = 1.15
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2 = 1.30
+ sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2 = 1.30
+ sky130_fd_pr__rf_pfet_01v8__aw_rd_mult = 1.0
+ sky130_fd_pr__rf_pfet_01v8__aw_rs_mult = 1.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_0 = -0.026318
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_0 = -0.00026051
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_0 = 0.036371
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_0 = 9011.9
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_0 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_1 = -0.0083086
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_1 = -0.00025544
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_1 = 0.043744
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_1 = -13691.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_1 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_2 = 0.00092097
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_2 = -0.00036227
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_2 = 0.025821
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_2 = -12946.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_2 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_3 = -0.023482
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_3 = -0.00065054
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_3 = 0.062883
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_3 = -10906.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_3 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_4 = -0.018913
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_4 = -0.00048132
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_4 = 0.054592
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_4 = -4787.1
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_4 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_5 = -0.016498
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_5 = -0.00040228
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_5 = 0.025581
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_5 = -7701.6
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_5 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_6 = -0.02415
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_6 = -0.0010764
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_6 = 0.088259
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_6 = -9692.8
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_7 = -0.00045958
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_7 = -12867.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_7 = -0.013677
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_7 = 0.054734
*
* sky130_fd_pr__rf_pfet_01v8_bM02, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM02__vth0_diff_8 = 0.03218
+ sky130_fd_pr__rf_pfet_01v8_bM02__u0_diff_8 = -0.00053308
+ sky130_fd_pr__rf_pfet_01v8_bM02__vsat_diff_8 = -16884.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ub_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM02__k2_diff_8 = -0.012368
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 000, W = 1.65, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_0 = -0.025153
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_0 = -0.00045786
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_0 = 0.049883
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_0 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_0 = 4304.4
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 001, W = 1.65, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_1 = -0.0081868
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_1 = -0.0003546
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_1 = 0.058034
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_1 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_1 = -1647.5
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 002, W = 1.65, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_2 = -0.00039936
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_2 = 0.0326
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_2 = -10830.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_2 = -0.00049705
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_2 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_2 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 003, W = 3.01, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_3 = -0.021287
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_3 = -0.00070687
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_3 = 0.061799
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_3 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_3 = -10201.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 004, W = 3.01, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_4 = -0.00073938
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_4 = 0.067454
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_4 = -10506.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_4 = -0.015399
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_4 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_4 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 005, W = 3.01, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_5 = 0.033162
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_5 = -0.00052171
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_5 = -14143.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_5 = -0.016662
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_5 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_5 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 006, W = 5.05, L = 0.15
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_6 = 0.091648
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_6 = -0.00096119
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_6 = -7280.9
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_6 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_6 = -0.023369
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 007, W = 5.05, L = 0.18
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_7 = -0.010709
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_7 = 0.059069
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_7 = -0.0007366
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_7 = -12730.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_7 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_7 = 0.0
*
* sky130_fd_pr__rf_pfet_01v8_bM04, Bin 008, W = 5.05, L = 0.25
* ------------------------------------------------
+ sky130_fd_pr__rf_pfet_01v8_bM04__rdsw_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__k2_diff_8 = -0.0113
+ sky130_fd_pr__rf_pfet_01v8_bM04__kt1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__nfactor_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ags_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__a0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__voff_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b0_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vth0_diff_8 = 0.044518
+ sky130_fd_pr__rf_pfet_01v8_bM04__u0_diff_8 = -0.00066793
+ sky130_fd_pr__rf_pfet_01v8_bM04__ua_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__vsat_diff_8 = -13679.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__b1_diff_8 = 0.0
+ sky130_fd_pr__rf_pfet_01v8_bM04__ub_diff_8 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__rf_pfet_01v8_b.pm3.spice"
