* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param
+ sky130_fd_pr__nfet_20v0__toxe_mult = 1.0
+ sky130_fd_pr__nfet_20v0__rshn_mult = 1.0
+ sky130_fd_pr__nfet_20v0__overlap_mult = 0.89805
+ sky130_fd_pr__nfet_20v0__ajunction_mult = 9.9505e-1
+ sky130_fd_pr__nfet_20v0__pjunction_mult = 1.0144
+ sky130_fd_pr__nfet_20v0__lint_diff = 0.0
+ sky130_fd_pr__nfet_20v0__wint_diff = 0.0
+ sky130_fd_pr__nfet_20v0__dlc_diff = 0.0
+ sky130_fd_pr__nfet_20v0__dwc_diff = 0.0
*
* sky130_fd_pr__nfet_20v0, Bin 000, W = 30.0u, L = 1.0u
* -----------------------------------
.param
+ sky130_fd_pr__nfet_20v0__rdrift_mult = 9.6982e-1
+ sky130_fd_pr__nfet_20v0__hvvsat_mult = 9.2197e-1
+ sky130_fd_pr__nfet_20v0__vth0_diff = 3.4824e-2
+ sky130_fd_pr__nfet_20v0__k2_diff = -2.7400e-2
*
* sky130_fd_pr__nfet_20v0_iso, Bin 000, W = 30.0u, L = 1.0u
* --------------------------------------
.param
+ sky130_fd_pr__nfet_20v0_iso__rdrift_mult = 9.1661e-1
+ sky130_fd_pr__nfet_20v0_iso__hvvsat_mult = 8.5177e-1
+ sky130_fd_pr__nfet_20v0_iso__vth0_diff = -1.2392e-3
+ sky130_fd_pr__nfet_20v0_iso__k2_diff = -1.9873e-2
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_20v0__subcircuit.pm3.spice"
*.include "sky130_fd_pr_models/nfet_20v0_iso/sky130_fd_pr__nfet_20v0_iso__subcircuit.pm3.spice"
*.include "sky130_fd_pr_models/nfet_20v0_zvt/sky130_fd_pr__nfet_20v0_zvt__tt_discrete.corner.spice"
.include "sky130_fd_pr_models/sky130_fd_pr__nfet_20v0_iso__subcircuit.pm3.spice"
.include "sky130_fd_pr_models/sky130_fd_pr__nfet_20v0_zvt__tt_discrete.corner.spice"
