* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.include "sky130_fd_pr_models/parasitics/sky130_fd_pr__model__parasitic__diode_pw2dn.model.spice"
.include "sky130_fd_pr_models/parasitics/sky130_fd_pr__model__parasitic__diode_pw2dn_noresistor.model.spice"
.include "sky130_fd_pr_models/parasitics/sky130_fd_pr__model__parasitic__rf_diode_pw2dn.model.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__esd_rf_diode_pw2nd_11v0_100__parasitic__diode_pw2dn.model.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__esd_rf_diode_pw2nd_11v0_200__parasitic__diode_pw2dn.model.spice"
.include "sky130_fd_pr_models/cells/sky130_fd_pr__esd_rf_diode_pw2nd_11v0_300__parasitic__diode_pw2dn.model.spice"
