* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* statistics {
* 	mismatch {
*     	}
*         process {
* 		vary sky130_fd_pr__res_xhigh_po__var_mult dist=gauss std=0.025
* 		vary sky130_fd_pr__res_high_po__var       dist=gauss std=0.025
*         }
* }
.subckt  sky130_fd_pr__model__parasitic__res_po r0 r1 sub
+ w=1u l=1u
*c0 r0 sub  c = {((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_1_1*1e-6)/2}    ; _option_scale_
*c1 r1 sub  c = {((l+2*2.08)*w*crpf_precision*1e-12+2*(l+2*2.08+w)*crpfsw_precision_1_1*1e-6)/2}    ; _option_scale_
c0 r0 sub  c = {((l+2*2.08e-6)*w*crpf_precision+2*((l+2*2.08e-6)+w)*crpfsw_precision_1_1)/2}
c1 r1 sub  c = {((l+2*2.08e-6)*w*crpf_precision+2*((l+2*2.08e-6)+w)*crpfsw_precision_1_1)/2}
.ends sky130_fd_pr__model__parasitic__res_po
