* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_01v8 d g s b
+ 
.param  l = 1u w = 1u ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 nf = 1.0
msky130_fd_pr__pfet_01v8 d g s b sky130_fd_pr__pfet_01v8__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
.model sky130_fd_pr__pfet_01v8__model.0 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.255e-06 wmax = 1.265e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0652+sky130_fd_pr__pfet_01v8__vth0_diff_0+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3152469
+ k2 = {-0.27798063+sky130_fd_pr__pfet_01v8__k2_diff_0}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {68611+sky130_fd_pr__pfet_01v8__vsat_diff_0}
+ ua = {-2.4423e-009+sky130_fd_pr__pfet_01v8__ua_diff_0}
+ ub = {2.0699352e-018+sky130_fd_pr__pfet_01v8__ub_diff_0}
+ uc = 1.6133739e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_0}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0025134+sky130_fd_pr__pfet_01v8__u0_diff_0}
+ a0 = {0.91285081+sky130_fd_pr__pfet_01v8__a0_diff_0}
+ keta = {-0.020464881+sky130_fd_pr__pfet_01v8__keta_diff_0}
+ a1 = 0.0
+ a2 = 0.87366558
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_0}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_0}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_0}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.25076476+sky130_fd_pr__pfet_01v8__voff_diff_0+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_0+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_0}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.21064695+sky130_fd_pr__pfet_01v8__eta0_diff_0}
+ etab = -0.014728557
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.61630162+sky130_fd_pr__pfet_01v8__pclm_diff_0}
+ pdiblc1 = 0.14215108
+ pdiblc2 = 0.0026509038
+ pdiblcb = -0.15188768
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.1788025e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.9381315
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_0}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_0}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {4.0078966e-010+sky130_fd_pr__pfet_01v8__agidl_diff_0}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_0}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_0}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_0}
+ kt2 = -0.12
+ at = 50942.0
+ ute = -0.21243
+ ua1 = 1.8303e-10
+ ub1 = 3.6891e-19
+ uc1 = 6.4484e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.1 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.675e-06 wmax = 1.685e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.02+sky130_fd_pr__pfet_01v8__vth0_diff_1+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3255051
+ k2 = {-0.28016116+sky130_fd_pr__pfet_01v8__k2_diff_1}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {59524+sky130_fd_pr__pfet_01v8__vsat_diff_1}
+ ua = {-2.4816e-009+sky130_fd_pr__pfet_01v8__ua_diff_1}
+ ub = {2.1055982e-018+sky130_fd_pr__pfet_01v8__ub_diff_1}
+ uc = 9.1597053e-14
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_1}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0024424+sky130_fd_pr__pfet_01v8__u0_diff_1}
+ a0 = {0.80890904+sky130_fd_pr__pfet_01v8__a0_diff_1}
+ keta = {0.027840733+sky130_fd_pr__pfet_01v8__keta_diff_1}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_1}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_1}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_1}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.27372667+sky130_fd_pr__pfet_01v8__voff_diff_1+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_1+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_1}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.3010182+sky130_fd_pr__pfet_01v8__eta0_diff_1}
+ etab = -0.035338434
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.47998966+sky130_fd_pr__pfet_01v8__pclm_diff_1}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.4222865e-5
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3226724e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.537679
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_1}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_1}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.8211658e-010+sky130_fd_pr__pfet_01v8__agidl_diff_1}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_1}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_1}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_1}
+ kt2 = -0.12
+ at = 39225.0
+ ute = -0.21243
+ ua1 = 1.6473e-10
+ ub1 = 3.6891e-19
+ uc1 = 6.4484e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.2 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.005+sky130_fd_pr__pfet_01v8__vth0_diff_2+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.45361058
+ k2 = {0.017567785+sky130_fd_pr__pfet_01v8__k2_diff_2}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {28810.641+sky130_fd_pr__pfet_01v8__vsat_diff_2}
+ ua = {-7.4785951e-010+sky130_fd_pr__pfet_01v8__ua_diff_2}
+ ub = {6.5707758e-019+sky130_fd_pr__pfet_01v8__ub_diff_2}
+ uc = -4.8679745e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_2}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0072271+sky130_fd_pr__pfet_01v8__u0_diff_2}
+ a0 = {0.63175+sky130_fd_pr__pfet_01v8__a0_diff_2}
+ keta = {-0.037840736+sky130_fd_pr__pfet_01v8__keta_diff_2}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {1.153125+sky130_fd_pr__pfet_01v8__ags_diff_2}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_2}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_2}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17660159+sky130_fd_pr__pfet_01v8__voff_diff_2+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_2+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_2}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_2}
+ etab = -0.007
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.37137649+sky130_fd_pr__pfet_01v8__pclm_diff_2}
+ pdiblc1 = 0.38223933
+ pdiblc2 = 0.000215
+ pdiblcb = -0.025
+ drout = 0.9112528
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.4098587e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.9010262
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_2}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_2}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_2}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_2}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_2}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.51384673+sky130_fd_pr__pfet_01v8__kt1_diff_2}
+ kt2 = -0.06387541
+ at = 22950.061
+ ute = -1.1934315
+ ua1 = -2.4046243e-10
+ ub1 = 4.7991978e-19
+ uc1 = 4.7436576e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.3 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0193+sky130_fd_pr__pfet_01v8__vth0_diff_3+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.46123612
+ k2 = {0.019412161+sky130_fd_pr__pfet_01v8__k2_diff_3}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {53437.5+sky130_fd_pr__pfet_01v8__vsat_diff_3}
+ ua = {-1.0211363e-009+sky130_fd_pr__pfet_01v8__ua_diff_3}
+ ub = {7.9306706e-019+sky130_fd_pr__pfet_01v8__ub_diff_3}
+ uc = -4.5032348e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_3}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.006259+sky130_fd_pr__pfet_01v8__u0_diff_3}
+ a0 = {1.1302+sky130_fd_pr__pfet_01v8__a0_diff_3}
+ keta = {-0.0048142243+sky130_fd_pr__pfet_01v8__keta_diff_3}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.37980837+sky130_fd_pr__pfet_01v8__ags_diff_3}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_3}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_3}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17603939+sky130_fd_pr__pfet_01v8__voff_diff_3+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5884088+sky130_fd_pr__pfet_01v8__nfactor_diff_3+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_3}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.0005+sky130_fd_pr__pfet_01v8__eta0_diff_3}
+ etab = -0.00050000149
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.35228743+sky130_fd_pr__pfet_01v8__pclm_diff_3}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3721337e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.048987e-12
+ alpha1 = -2.9238605e-15
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_3}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_3}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.4838246e-010+sky130_fd_pr__pfet_01v8__agidl_diff_3}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_3}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_3}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47097+sky130_fd_pr__pfet_01v8__kt1_diff_3}
+ kt2 = -0.045529
+ at = 7459.5
+ ute = -0.89505
+ ua1 = -1.5331e-10
+ ub1 = 7.4669e-19
+ uc1 = 6.1866e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.4 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.01+sky130_fd_pr__pfet_01v8__vth0_diff_4+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44975853
+ k2 = {0.023544581+sky130_fd_pr__pfet_01v8__k2_diff_4}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {42745.77+sky130_fd_pr__pfet_01v8__vsat_diff_4}
+ ua = {-8.2697914e-010+sky130_fd_pr__pfet_01v8__ua_diff_4}
+ ub = {6.6035544e-019+sky130_fd_pr__pfet_01v8__ub_diff_4}
+ uc = -5.4570621e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_4}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0068894+sky130_fd_pr__pfet_01v8__u0_diff_4}
+ a0 = {1.1794+sky130_fd_pr__pfet_01v8__a0_diff_4}
+ keta = {0.0032223923+sky130_fd_pr__pfet_01v8__keta_diff_4}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.29875546+sky130_fd_pr__pfet_01v8__ags_diff_4}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_4}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_4}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1748426+sky130_fd_pr__pfet_01v8__voff_diff_4+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_4+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_4}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_4}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.038003634+sky130_fd_pr__pfet_01v8__pclm_diff_4}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0010378863
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 7.9999998e+8
+ pscbe2 = 9.5028802e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_4}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_4}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.5747859e-010+sky130_fd_pr__pfet_01v8__agidl_diff_4}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_4}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_4}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.46128+sky130_fd_pr__pfet_01v8__kt1_diff_4}
+ kt2 = -0.026742
+ at = 55268.5
+ ute = -0.07
+ ua1 = 1.9196e-9
+ ub1 = -1.0155e-18
+ uc1 = -8.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.5 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.99608+sky130_fd_pr__pfet_01v8__vth0_diff_5+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.49177002
+ k2 = {0.012599753+sky130_fd_pr__pfet_01v8__k2_diff_5}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {55237.817+sky130_fd_pr__pfet_01v8__vsat_diff_5}
+ ua = {-1.3880621e-009+sky130_fd_pr__pfet_01v8__ua_diff_5}
+ ub = {1.048282e-018+sky130_fd_pr__pfet_01v8__ub_diff_5}
+ uc = -3.8916596e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_5}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0048205252+sky130_fd_pr__pfet_01v8__u0_diff_5}
+ a0 = {1.29386+sky130_fd_pr__pfet_01v8__a0_diff_5}
+ keta = {0.0066402373+sky130_fd_pr__pfet_01v8__keta_diff_5}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.20242817+sky130_fd_pr__pfet_01v8__ags_diff_5}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_5}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_5}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17895891+sky130_fd_pr__pfet_01v8__voff_diff_5+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4721938+sky130_fd_pr__pfet_01v8__nfactor_diff_5+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_5}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_5}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.0017402344+sky130_fd_pr__pfet_01v8__pclm_diff_5}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 7.9998529e+8
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_5}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_5}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.4670794e-010+sky130_fd_pr__pfet_01v8__agidl_diff_5}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_5}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_5}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.54561+sky130_fd_pr__pfet_01v8__kt1_diff_5}
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.6 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97755+sky130_fd_pr__pfet_01v8__vth0_diff_6+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.4974388
+ k2 = {-0.34240453+sky130_fd_pr__pfet_01v8__k2_diff_6}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {55335+sky130_fd_pr__pfet_01v8__vsat_diff_6}
+ ua = {-2.5669e-009+sky130_fd_pr__pfet_01v8__ua_diff_6}
+ ub = {2.1902542e-018+sky130_fd_pr__pfet_01v8__ub_diff_6}
+ uc = 2.3206046e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_6}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0020949+sky130_fd_pr__pfet_01v8__u0_diff_6}
+ a0 = {0.72595373+sky130_fd_pr__pfet_01v8__a0_diff_6}
+ keta = {-0.0003767501+sky130_fd_pr__pfet_01v8__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_6}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_6}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28041511+sky130_fd_pr__pfet_01v8__voff_diff_6+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.892779+sky130_fd_pr__pfet_01v8__nfactor_diff_6+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_6}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.34230525+sky130_fd_pr__pfet_01v8__eta0_diff_6}
+ etab = -1.1566507e-13
+ dsub = 0.26628854
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.45374464+sky130_fd_pr__pfet_01v8__pclm_diff_6}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.4414063e-5
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3761341e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.2512308
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.1989212e-010+sky130_fd_pr__pfet_01v8__agidl_diff_6}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_6}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_6}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_6}
+ kt2 = -0.12
+ at = 21109.0
+ ute = -0.21243
+ ua1 = 1.0762e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.7 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.95759+sky130_fd_pr__pfet_01v8__vth0_diff_7+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.1286524
+ k2 = {-0.20642701+sky130_fd_pr__pfet_01v8__k2_diff_7}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {81677+sky130_fd_pr__pfet_01v8__vsat_diff_7}
+ ua = {-2.3466042e-009+sky130_fd_pr__pfet_01v8__ua_diff_7}
+ ub = {1.9914931e-018+sky130_fd_pr__pfet_01v8__ub_diff_7}
+ uc = 2.2913949e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_7}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0027565+sky130_fd_pr__pfet_01v8__u0_diff_7}
+ a0 = {1.087+sky130_fd_pr__pfet_01v8__a0_diff_7}
+ keta = {0.027122826+sky130_fd_pr__pfet_01v8__keta_diff_7}
+ a1 = 0.0
+ a2 = 0.68678659
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_7}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_7}
+ b1 = {2.1073424e-024+sky130_fd_pr__pfet_01v8__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.24161658+sky130_fd_pr__pfet_01v8__voff_diff_7+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_7+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_7}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.21136947+sky130_fd_pr__pfet_01v8__eta0_diff_7}
+ etab = -0.031554764
+ dsub = 0.26948731
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62205899+sky130_fd_pr__pfet_01v8__pclm_diff_7}
+ pdiblc1 = 0.15224245
+ pdiblc2 = 0.0023148811
+ pdiblcb = -0.075
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3883381e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.7923713
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_7}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_7}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_7}
+ bgidl = {1.0029534e009+sky130_fd_pr__pfet_01v8__bgidl_diff_7}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_7}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.63808+sky130_fd_pr__pfet_01v8__kt1_diff_7}
+ kt2 = -0.12
+ at = 59144.0
+ ute = -0.21616
+ ua1 = 1.505e-10
+ ub1 = 4.39e-19
+ uc1 = 9.4135e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.8 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.99068+sky130_fd_pr__pfet_01v8__vth0_diff_8+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 0.58024567
+ k2 = {-0.012344333+sky130_fd_pr__pfet_01v8__k2_diff_8}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {123990.79+sky130_fd_pr__pfet_01v8__vsat_diff_8}
+ ua = {-1.5758775e-009+sky130_fd_pr__pfet_01v8__ua_diff_8}
+ ub = {1.3921314e-018+sky130_fd_pr__pfet_01v8__ub_diff_8}
+ uc = 5.5432313e-14
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_8}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0054984+sky130_fd_pr__pfet_01v8__u0_diff_8}
+ a0 = {0.81211+sky130_fd_pr__pfet_01v8__a0_diff_8}
+ keta = {-0.0099696456+sky130_fd_pr__pfet_01v8__keta_diff_8}
+ a1 = 0.0
+ a2 = 0.52372326
+ ags = {0.42180356+sky130_fd_pr__pfet_01v8__ags_diff_8}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_8}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_8}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.21482801+sky130_fd_pr__pfet_01v8__voff_diff_8+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_8+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_8}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_8}
+ etab = -6.25e-5
+ dsub = 0.62800029
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63715328+sky130_fd_pr__pfet_01v8__pclm_diff_8}
+ pdiblc1 = 0.46195031
+ pdiblc2 = 0.011067434
+ pdiblcb = -0.225
+ drout = 0.43167959
+ pscbe1 = 7.9992886e+8
+ pscbe2 = 9.2096719e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.2931629
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_8}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_8}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_8}
+ bgidl = {1.2773568e009+sky130_fd_pr__pfet_01v8__bgidl_diff_8}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_8}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.51207+sky130_fd_pr__pfet_01v8__kt1_diff_8}
+ kt2 = -0.017592
+ at = 66556.0
+ ute = -0.18527
+ ua1 = 4.0254e-10
+ ub1 = 4.39e-19
+ uc1 = 5.7234e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.9 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1+sky130_fd_pr__pfet_01v8__vth0_diff_9+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.50911445
+ k2 = {0.0041427676+sky130_fd_pr__pfet_01v8__k2_diff_9}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {74041+sky130_fd_pr__pfet_01v8__vsat_diff_9}
+ ua = {-1.1297907e-009+sky130_fd_pr__pfet_01v8__ua_diff_9}
+ ub = {9.744598e-019+sky130_fd_pr__pfet_01v8__ub_diff_9}
+ uc = -2.1796978e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_9}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0062005+sky130_fd_pr__pfet_01v8__u0_diff_9}
+ a0 = {1.1353+sky130_fd_pr__pfet_01v8__a0_diff_9}
+ keta = {-0.033356713+sky130_fd_pr__pfet_01v8__keta_diff_9}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {1.3126648+sky130_fd_pr__pfet_01v8__ags_diff_9}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_9}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_9}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1859804+sky130_fd_pr__pfet_01v8__voff_diff_9+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_9+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_9}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_9}
+ etab = -6.25e-6
+ dsub = 0.31741848
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62622696+sky130_fd_pr__pfet_01v8__pclm_diff_9}
+ pdiblc1 = 0.15515165
+ pdiblc2 = 0.00053219225
+ pdiblcb = -0.025
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.317151e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.0318843
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_9}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_9}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.7836505e-010+sky130_fd_pr__pfet_01v8__agidl_diff_9}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_9}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_9}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.50846+sky130_fd_pr__pfet_01v8__kt1_diff_9}
+ kt2 = -0.055188
+ at = 65000.0
+ ute = -0.24063
+ ua1 = 5.5621e-10
+ ub1 = 5.5151e-19
+ uc1 = 2.432e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.10 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.995e-06 wmax = 2.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97864+sky130_fd_pr__pfet_01v8__vth0_diff_10+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.4657817
+ k2 = {-0.34178317+sky130_fd_pr__pfet_01v8__k2_diff_10}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {58358+sky130_fd_pr__pfet_01v8__vsat_diff_10}
+ ua = {-2.5888e-009+sky130_fd_pr__pfet_01v8__ua_diff_10}
+ ub = {2.2070427e-018+sky130_fd_pr__pfet_01v8__ub_diff_10}
+ uc = 1.0397944e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_10}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0021842+sky130_fd_pr__pfet_01v8__u0_diff_10}
+ a0 = {0.57015042+sky130_fd_pr__pfet_01v8__a0_diff_10}
+ keta = {-0.038910431+sky130_fd_pr__pfet_01v8__keta_diff_10}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {0.0640625+sky130_fd_pr__pfet_01v8__ags_diff_10}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_10}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_10}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.27300243+sky130_fd_pr__pfet_01v8__voff_diff_10+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_10+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_10}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.28103229+sky130_fd_pr__pfet_01v8__eta0_diff_10}
+ etab = -2.7452546e-151
+ dsub = 0.26029894
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.53574449+sky130_fd_pr__pfet_01v8__pclm_diff_10}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.0
+ pscbe1 = 7.8140327e+8
+ pscbe2 = 9.2985538e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.4455034
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_10}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_10}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.4770616e-010+sky130_fd_pr__pfet_01v8__agidl_diff_10}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_10}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_10}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_10}
+ kt2 = -0.12
+ at = 25889.0
+ ute = -0.21243
+ ua1 = 1.3508e-10
+ ub1 = 3.8367e-19
+ uc1 = 6.4484e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.11 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1+sky130_fd_pr__pfet_01v8__vth0_diff_11+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.48077988
+ k2 = {0.016877332+sky130_fd_pr__pfet_01v8__k2_diff_11}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {52076.876+sky130_fd_pr__pfet_01v8__vsat_diff_11}
+ ua = {-1.3191618e-009+sky130_fd_pr__pfet_01v8__ua_diff_11}
+ ub = {9.9701215e-019+sky130_fd_pr__pfet_01v8__ub_diff_11}
+ uc = -3.009708e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_11}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.005252+sky130_fd_pr__pfet_01v8__u0_diff_11}
+ a0 = {1.139+sky130_fd_pr__pfet_01v8__a0_diff_11}
+ keta = {-0.0079115309+sky130_fd_pr__pfet_01v8__keta_diff_11}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.57328989+sky130_fd_pr__pfet_01v8__ags_diff_11}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_11}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_11}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19564023+sky130_fd_pr__pfet_01v8__voff_diff_11+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3744146+sky130_fd_pr__pfet_01v8__nfactor_diff_11+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_11}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_11}
+ etab = -22.773578
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62700535+sky130_fd_pr__pfet_01v8__pclm_diff_11}
+ pdiblc1 = 0.37610116
+ pdiblc2 = 0.00043
+ pdiblcb = -0.00077709656
+ drout = 0.75941084
+ pscbe1 = 8.0e+8
+ pscbe2 = 7.3674496e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.8770833
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_11}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_11}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_11}
+ bgidl = {1.1984227e009+sky130_fd_pr__pfet_01v8__bgidl_diff_11}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_11}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.44959+sky130_fd_pr__pfet_01v8__kt1_diff_11}
+ kt2 = -0.050195
+ at = 64793.0
+ ute = -0.40685
+ ua1 = 2.5217e-10
+ ub1 = 5.1252e-19
+ uc1 = 9.446e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.12 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0251+sky130_fd_pr__pfet_01v8__vth0_diff_12+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.51320198
+ k2 = {-0.0022346833+sky130_fd_pr__pfet_01v8__k2_diff_12}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {24613.898+sky130_fd_pr__pfet_01v8__vsat_diff_12}
+ ua = {-7.9601337e-010+sky130_fd_pr__pfet_01v8__ua_diff_12}
+ ub = {6.5199713e-019+sky130_fd_pr__pfet_01v8__ub_diff_12}
+ uc = -6.4508638e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_12}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0071794+sky130_fd_pr__pfet_01v8__u0_diff_12}
+ a0 = {1.0021+sky130_fd_pr__pfet_01v8__a0_diff_12}
+ keta = {-0.021786634+sky130_fd_pr__pfet_01v8__keta_diff_12}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.53430225+sky130_fd_pr__pfet_01v8__ags_diff_12}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_12}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_12}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1918163+sky130_fd_pr__pfet_01v8__voff_diff_12+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5680269+sky130_fd_pr__pfet_01v8__nfactor_diff_12+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_12}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_12}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.41578123+sky130_fd_pr__pfet_01v8__pclm_diff_12}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0013376645
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.0332673e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0432903e-11
+ alpha1 = 1.0e-10
+ beta0 = 6.5167702
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_12}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_12}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.5891284e-010+sky130_fd_pr__pfet_01v8__agidl_diff_12}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_12}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_12}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47463+sky130_fd_pr__pfet_01v8__kt1_diff_12}
+ kt2 = -0.056201
+ at = 27226.0
+ ute = -1.0471
+ ua1 = -1.7587e-10
+ ub1 = 6.1469e-19
+ uc1 = 1.0103e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.13 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0425+sky130_fd_pr__pfet_01v8__vth0_diff_13+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.45544295
+ k2 = {0.017209681+sky130_fd_pr__pfet_01v8__k2_diff_13}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {29822.135+sky130_fd_pr__pfet_01v8__vsat_diff_13}
+ ua = {-2.8340104e-010+sky130_fd_pr__pfet_01v8__ua_diff_13}
+ ub = {3.9493106e-019+sky130_fd_pr__pfet_01v8__ub_diff_13}
+ uc = -8.5236227e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_13}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0095057+sky130_fd_pr__pfet_01v8__u0_diff_13}
+ a0 = {1.1338+sky130_fd_pr__pfet_01v8__a0_diff_13}
+ keta = {-0.0096897358+sky130_fd_pr__pfet_01v8__keta_diff_13}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.31273428+sky130_fd_pr__pfet_01v8__ags_diff_13}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_13}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_13}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20325421+sky130_fd_pr__pfet_01v8__voff_diff_13+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6422165+sky130_fd_pr__pfet_01v8__nfactor_diff_13+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_13}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_13}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.4127159+sky130_fd_pr__pfet_01v8__pclm_diff_13}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.5112332e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.4560427e-11
+ alpha1 = 8.8540421e-13
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_13}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_13}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.3573869e-010+sky130_fd_pr__pfet_01v8__agidl_diff_13}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_13}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_13}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.45286769+sky130_fd_pr__pfet_01v8__kt1_diff_13}
+ kt2 = -0.051427601
+ at = 46321.73
+ ute = -0.15559115
+ ua1 = 2.1813426e-9
+ ub1 = -9.2319056e-19
+ uc1 = -1.3034169e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.14 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0502+sky130_fd_pr__pfet_01v8__vth0_diff_14+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = {0.029470664+sky130_fd_pr__pfet_01v8__k2_diff_14}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {53438+sky130_fd_pr__pfet_01v8__vsat_diff_14}
+ ua = {-1.8971577e-010+sky130_fd_pr__pfet_01v8__ua_diff_14}
+ ub = {3.1380962e-019+sky130_fd_pr__pfet_01v8__ub_diff_14}
+ uc = -9.8608028e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_14}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0096116+sky130_fd_pr__pfet_01v8__u0_diff_14}
+ a0 = {1.1296+sky130_fd_pr__pfet_01v8__a0_diff_14}
+ keta = {4.9707517e-006+sky130_fd_pr__pfet_01v8__keta_diff_14}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.16627013+sky130_fd_pr__pfet_01v8__ags_diff_14}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_14}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_14}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.21413558+sky130_fd_pr__pfet_01v8__voff_diff_14+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.706221+sky130_fd_pr__pfet_01v8__nfactor_diff_14+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_14}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_14}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.14877095+sky130_fd_pr__pfet_01v8__pclm_diff_14}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.5712828e+8
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_14}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_14}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_14}
+ bgidl = {1.3525405e009+sky130_fd_pr__pfet_01v8__bgidl_diff_14}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_14}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.4443203+sky130_fd_pr__pfet_01v8__kt1_diff_14}
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.15 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.018+sky130_fd_pr__pfet_01v8__vth0_diff_15+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3168639
+ k2 = {-0.28483489+sky130_fd_pr__pfet_01v8__k2_diff_15}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {62767+sky130_fd_pr__pfet_01v8__vsat_diff_15}
+ ua = {-2.4824e-009+sky130_fd_pr__pfet_01v8__ua_diff_15}
+ ub = {2.1281765e-018+sky130_fd_pr__pfet_01v8__ub_diff_15}
+ uc = 1.970052e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_15}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0026317+sky130_fd_pr__pfet_01v8__u0_diff_15}
+ a0 = {0.84981148+sky130_fd_pr__pfet_01v8__a0_diff_15}
+ keta = {0.014244979+sky130_fd_pr__pfet_01v8__keta_diff_15}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_15}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_15}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_15}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.29628465+sky130_fd_pr__pfet_01v8__voff_diff_15+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_15+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_15}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.33076312+sky130_fd_pr__pfet_01v8__eta0_diff_15}
+ etab = -0.01389211
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.4433904+sky130_fd_pr__pfet_01v8__pclm_diff_15}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -4.8637071e-5
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.5586458e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.3823117
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_15}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_15}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.7158891e-010+sky130_fd_pr__pfet_01v8__agidl_diff_15}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_15}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_15}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.695+sky130_fd_pr__pfet_01v8__kt1_diff_15}
+ kt2 = -0.12196
+ at = 38000.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.16 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.004+sky130_fd_pr__pfet_01v8__vth0_diff_16+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.0376715
+ k2 = {-0.17335648+sky130_fd_pr__pfet_01v8__k2_diff_16}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {88456+sky130_fd_pr__pfet_01v8__vsat_diff_16}
+ ua = {-2.2421727e-009+sky130_fd_pr__pfet_01v8__ua_diff_16}
+ ub = {1.8536584e-018+sky130_fd_pr__pfet_01v8__ub_diff_16}
+ uc = 2.5234343e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_16}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0029971+sky130_fd_pr__pfet_01v8__u0_diff_16}
+ a0 = {0.89088+sky130_fd_pr__pfet_01v8__a0_diff_16}
+ keta = {0.023895141+sky130_fd_pr__pfet_01v8__keta_diff_16}
+ a1 = 0.0
+ a2 = 0.67187683
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_16}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_16}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_16}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22630768+sky130_fd_pr__pfet_01v8__voff_diff_16+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.7534082+sky130_fd_pr__pfet_01v8__nfactor_diff_16+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_16}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.18201237+sky130_fd_pr__pfet_01v8__eta0_diff_16}
+ etab = -0.078353952
+ dsub = 0.27170577
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63088962+sky130_fd_pr__pfet_01v8__pclm_diff_16}
+ pdiblc1 = 0.18080115
+ pdiblc2 = 0.0040267418
+ pdiblcb = -0.0001934424
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.4769552e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.580652
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_16}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_16}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.0157032e-010+sky130_fd_pr__pfet_01v8__agidl_diff_16}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_16}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_16}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.598+sky130_fd_pr__pfet_01v8__kt1_diff_16}
+ kt2 = -0.12196
+ at = 68317.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.17 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.964+sky130_fd_pr__pfet_01v8__vth0_diff_17+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 0.77076332
+ k2 = {-0.082949567+sky130_fd_pr__pfet_01v8__k2_diff_17}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {77620+sky130_fd_pr__pfet_01v8__vsat_diff_17}
+ ua = {-1.9102726e-009+sky130_fd_pr__pfet_01v8__ua_diff_17}
+ ub = {1.5401215e-018+sky130_fd_pr__pfet_01v8__ub_diff_17}
+ uc = -6.4335368e-12
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_17}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0041176+sky130_fd_pr__pfet_01v8__u0_diff_17}
+ a0 = {0.50091+sky130_fd_pr__pfet_01v8__a0_diff_17}
+ keta = {-0.077084505+sky130_fd_pr__pfet_01v8__keta_diff_17}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.90459965+sky130_fd_pr__pfet_01v8__ags_diff_17}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_17}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_17}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20537164+sky130_fd_pr__pfet_01v8__voff_diff_17+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.8793354+sky130_fd_pr__pfet_01v8__nfactor_diff_17+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_17}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.29288956+sky130_fd_pr__pfet_01v8__eta0_diff_17}
+ etab = -5.0000128e-5
+ dsub = 0.5018771
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.84907102+sky130_fd_pr__pfet_01v8__pclm_diff_17}
+ pdiblc1 = 0.38718759
+ pdiblc2 = 0.0077688684
+ pdiblcb = -0.12475545
+ drout = 0.58591194
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.2265127e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.9226154
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_17}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_17}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.5628906e-009+sky130_fd_pr__pfet_01v8__agidl_diff_17}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_17}
+ cgidl = {60.778499+sky130_fd_pr__pfet_01v8__cgidl_diff_17}
+ egidl = 1.3658824
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.53419+sky130_fd_pr__pfet_01v8__kt1_diff_17}
+ kt2 = -0.060854
+ at = 56209.0
+ ute = -0.3
+ ua1 = 2.0193e-10
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.18 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.992+sky130_fd_pr__pfet_01v8__vth0_diff_18+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.45068637
+ k2 = {0.032260684+sky130_fd_pr__pfet_01v8__k2_diff_18}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {73912+sky130_fd_pr__pfet_01v8__vsat_diff_18}
+ ua = {-1.2118425e-009+sky130_fd_pr__pfet_01v8__ua_diff_18}
+ ub = {1.0568551e-018+sky130_fd_pr__pfet_01v8__ub_diff_18}
+ uc = -7.1566623e-12
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_18}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.006132+sky130_fd_pr__pfet_01v8__u0_diff_18}
+ a0 = {1.0051+sky130_fd_pr__pfet_01v8__a0_diff_18}
+ keta = {-0.012396657+sky130_fd_pr__pfet_01v8__keta_diff_18}
+ a1 = 0.0
+ a2 = 0.84119211
+ ags = {1.0025754+sky130_fd_pr__pfet_01v8__ags_diff_18}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_18}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_18}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19696087+sky130_fd_pr__pfet_01v8__voff_diff_18+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3845847+sky130_fd_pr__pfet_01v8__nfactor_diff_18+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_18}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_18}
+ etab = -0.00046590341
+ dsub = 0.28932681
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62284281+sky130_fd_pr__pfet_01v8__pclm_diff_18}
+ pdiblc1 = 0.18912731
+ pdiblc2 = 0.00058741392
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3232486e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.3861845
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_18}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_18}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.0755899e-010+sky130_fd_pr__pfet_01v8__agidl_diff_18}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_18}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_18}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.50846+sky130_fd_pr__pfet_01v8__kt1_diff_18}
+ kt2 = -0.055188
+ at = 73880.0
+ ute = -0.31763
+ ua1 = 5.5621e-10
+ ub1 = 4.1736e-19
+ uc1 = 2.432e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.19 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0354+sky130_fd_pr__pfet_01v8__vth0_diff_19+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.51518623
+ k2 = {-0.0012746592+sky130_fd_pr__pfet_01v8__k2_diff_19}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {27963.813+sky130_fd_pr__pfet_01v8__vsat_diff_19}
+ ua = {-1.122802e-009+sky130_fd_pr__pfet_01v8__ua_diff_19}
+ ub = {9.9211788e-019+sky130_fd_pr__pfet_01v8__ub_diff_19}
+ uc = -3.022645e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_19}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0068302+sky130_fd_pr__pfet_01v8__u0_diff_19}
+ a0 = {0.73977+sky130_fd_pr__pfet_01v8__a0_diff_19}
+ keta = {-0.052199769+sky130_fd_pr__pfet_01v8__keta_diff_19}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {1.1223202+sky130_fd_pr__pfet_01v8__ags_diff_19}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_19}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_19}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19282254+sky130_fd_pr__pfet_01v8__voff_diff_19+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.803914+sky130_fd_pr__pfet_01v8__nfactor_diff_19+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_19}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_19}
+ etab = -0.0012500664
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.42072955+sky130_fd_pr__pfet_01v8__pclm_diff_19}
+ pdiblc1 = 0.38126049
+ pdiblc2 = 0.00043
+ pdiblcb = -0.00076262347
+ drout = 0.81189156
+ pscbe1 = 8.0e+8
+ pscbe2 = 7.2098721e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.9305788
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_19}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_19}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_19}
+ bgidl = {1.1834062e009+sky130_fd_pr__pfet_01v8__bgidl_diff_19}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_19}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47401239+sky130_fd_pr__pfet_01v8__kt1_diff_19}
+ kt2 = -0.047712156
+ at = 25416.096
+ ute = -0.23992986
+ ua1 = 1.9047573e-9
+ ub1 = -1.2373089e-18
+ uc1 = -1.1188284e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.20 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0434+sky130_fd_pr__pfet_01v8__vth0_diff_20+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.441928
+ k2 = {0.028912751+sky130_fd_pr__pfet_01v8__k2_diff_20}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {53437.5+sky130_fd_pr__pfet_01v8__vsat_diff_20}
+ ua = {-9.8137786e-010+sky130_fd_pr__pfet_01v8__ua_diff_20}
+ ub = {9.0965495e-019+sky130_fd_pr__pfet_01v8__ub_diff_20}
+ uc = -3.4413404e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_20}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0073345+sky130_fd_pr__pfet_01v8__u0_diff_20}
+ a0 = {1.1942+sky130_fd_pr__pfet_01v8__a0_diff_20}
+ keta = {-0.016745386+sky130_fd_pr__pfet_01v8__keta_diff_20}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.42664895+sky130_fd_pr__pfet_01v8__ags_diff_20}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_20}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_20}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20413517+sky130_fd_pr__pfet_01v8__voff_diff_20+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.313002+sky130_fd_pr__pfet_01v8__nfactor_diff_20+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_20}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.00050000191+sky130_fd_pr__pfet_01v8__eta0_diff_20}
+ etab = -0.00050000042
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.6390771+sky130_fd_pr__pfet_01v8__pclm_diff_20}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.8845095e+8
+ pscbe2 = 9.4549435e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.2326697
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_20}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_20}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_20}
+ bgidl = {1.3452252e009+sky130_fd_pr__pfet_01v8__bgidl_diff_20}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_20}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.46529126+sky130_fd_pr__pfet_01v8__kt1_diff_20}
+ kt2 = -0.044800084
+ at = 79543.736
+ ute = -0.29475285
+ ua1 = 1.4994695e-9
+ ub1 = -5.4876923e-19
+ uc1 = 1.1407361e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.21 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0554+sky130_fd_pr__pfet_01v8__vth0_diff_21+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.41493399
+ k2 = {0.038381535+sky130_fd_pr__pfet_01v8__k2_diff_21}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {56763.737+sky130_fd_pr__pfet_01v8__vsat_diff_21}
+ ua = {-3.9589575e-010+sky130_fd_pr__pfet_01v8__ua_diff_21}
+ ub = {5.1890668e-019+sky130_fd_pr__pfet_01v8__ub_diff_21}
+ uc = -6.119559e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_21}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0094763+sky130_fd_pr__pfet_01v8__u0_diff_21}
+ a0 = {1.1906+sky130_fd_pr__pfet_01v8__a0_diff_21}
+ keta = {-0.010442146+sky130_fd_pr__pfet_01v8__keta_diff_21}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.30079431+sky130_fd_pr__pfet_01v8__ags_diff_21}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_21}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_21}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20758432+sky130_fd_pr__pfet_01v8__voff_diff_21+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4973257+sky130_fd_pr__pfet_01v8__nfactor_diff_21+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_21}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_21}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.44022027+sky130_fd_pr__pfet_01v8__pclm_diff_21}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0001075
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.4653461e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.6700366
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_21}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_21}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_21}
+ bgidl = {1.4866338e009+sky130_fd_pr__pfet_01v8__bgidl_diff_21}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_21}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.46286769+sky130_fd_pr__pfet_01v8__kt1_diff_21}
+ kt2 = -0.051427601
+ at = 094321.73
+ ute = -0.20559115
+ ua1 = 2.1813426e-9
+ ub1 = -9.2319056e-19
+ uc1 = -1.3034169e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.22 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0559+sky130_fd_pr__pfet_01v8__vth0_diff_22+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43056354
+ k2 = {0.033552779+sky130_fd_pr__pfet_01v8__k2_diff_22}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {160312.5+sky130_fd_pr__pfet_01v8__vsat_diff_22}
+ ua = {-5.5284971e-010+sky130_fd_pr__pfet_01v8__ua_diff_22}
+ ub = {5.7443771e-019+sky130_fd_pr__pfet_01v8__ub_diff_22}
+ uc = -6.3227866e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_22}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0085639+sky130_fd_pr__pfet_01v8__u0_diff_22}
+ a0 = {1.2059+sky130_fd_pr__pfet_01v8__a0_diff_22}
+ keta = {-0.0048615622+sky130_fd_pr__pfet_01v8__keta_diff_22}
+ a1 = 0.0
+ a2 = 0.90977388
+ ags = {0.21791559+sky130_fd_pr__pfet_01v8__ags_diff_22}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_22}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_22}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.21105937+sky130_fd_pr__pfet_01v8__voff_diff_22+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5008954+sky130_fd_pr__pfet_01v8__nfactor_diff_22+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_22}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_22}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.22728372+sky130_fd_pr__pfet_01v8__pclm_diff_22}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00016870007
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.077064e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.3511639
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_22}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_22}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_22}
+ bgidl = {1.5424014e009+sky130_fd_pr__pfet_01v8__bgidl_diff_22}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_22}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.43605364+sky130_fd_pr__pfet_01v8__kt1_diff_22}
+ kt2 = -0.050535666
+ at = 90000.0
+ ute = -0.16471211
+ ua1 = 1.9593569e-9
+ ub1 = -7.5242716e-19
+ uc1 = 1.1193066e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.23 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0213+sky130_fd_pr__pfet_01v8__vth0_diff_23+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.292041
+ k2 = {-0.27943118+sky130_fd_pr__pfet_01v8__k2_diff_23}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {68644+sky130_fd_pr__pfet_01v8__vsat_diff_23}
+ ua = {-2.5207e-009+sky130_fd_pr__pfet_01v8__ua_diff_23}
+ ub = {2.1497621e-018+sky130_fd_pr__pfet_01v8__ub_diff_23}
+ uc = 1.3933536e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_23}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0026411+sky130_fd_pr__pfet_01v8__u0_diff_23}
+ a0 = {0.95628558+sky130_fd_pr__pfet_01v8__a0_diff_23}
+ keta = {-0.0098450238+sky130_fd_pr__pfet_01v8__keta_diff_23}
+ a1 = 0.0
+ a2 = 0.83110554
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_23}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_23}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_23}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26814403+sky130_fd_pr__pfet_01v8__voff_diff_23+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_23+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_23}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.29347494+sky130_fd_pr__pfet_01v8__eta0_diff_23}
+ etab = -0.014445067
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.46055509+sky130_fd_pr__pfet_01v8__pclm_diff_23}
+ pdiblc1 = 0.019500056
+ pdiblc2 = 0.0014727467
+ pdiblcb = -0.075
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3135595e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.6984199
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_23}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_23}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.3920965e-010+sky130_fd_pr__pfet_01v8__agidl_diff_23}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_23}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_23}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.693+sky130_fd_pr__pfet_01v8__kt1_diff_23}
+ kt2 = -0.12196
+ at = 38000.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.24 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.004+sky130_fd_pr__pfet_01v8__vth0_diff_24+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.035054
+ k2 = {-0.17495984+sky130_fd_pr__pfet_01v8__k2_diff_24}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {77466+sky130_fd_pr__pfet_01v8__vsat_diff_24}
+ ua = {-2.2596593e-009+sky130_fd_pr__pfet_01v8__ua_diff_24}
+ ub = {1.8740807e-018+sky130_fd_pr__pfet_01v8__ub_diff_24}
+ uc = 2.1939953e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_24}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0032489+sky130_fd_pr__pfet_01v8__u0_diff_24}
+ a0 = {0.51935+sky130_fd_pr__pfet_01v8__a0_diff_24}
+ keta = {-0.049156996+sky130_fd_pr__pfet_01v8__keta_diff_24}
+ a1 = 0.0
+ a2 = 0.76127491
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_24}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_24}
+ b1 = {2.1073424e-024+sky130_fd_pr__pfet_01v8__b1_diff_24}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.24011109+sky130_fd_pr__pfet_01v8__voff_diff_24+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_24+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_24}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.19769484+sky130_fd_pr__pfet_01v8__eta0_diff_24}
+ etab = -0.055771336
+ dsub = 0.30311035
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63770979+sky130_fd_pr__pfet_01v8__pclm_diff_24}
+ pdiblc1 = 0.19075739
+ pdiblc2 = 0.004218602
+ pdiblcb = -0.075
+ drout = 0.91135477
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3641435e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.5831969
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_24}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_24}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_24}
+ bgidl = {1.0931445e009+sky130_fd_pr__pfet_01v8__bgidl_diff_24}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_24}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.568+sky130_fd_pr__pfet_01v8__kt1_diff_24}
+ kt2 = -0.1183
+ at = 53240.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 1.5093e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.25 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.96902+sky130_fd_pr__pfet_01v8__vth0_diff_25+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 0.82329436
+ k2 = {-0.099569738+sky130_fd_pr__pfet_01v8__k2_diff_25}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {76519+sky130_fd_pr__pfet_01v8__vsat_diff_25}
+ ua = {-2.045889e-009+sky130_fd_pr__pfet_01v8__ua_diff_25}
+ ub = {1.6358053e-018+sky130_fd_pr__pfet_01v8__ub_diff_25}
+ uc = 1.1896412e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_25}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0037126+sky130_fd_pr__pfet_01v8__u0_diff_25}
+ a0 = {0.66876525+sky130_fd_pr__pfet_01v8__a0_diff_25}
+ keta = {-0.10104013+sky130_fd_pr__pfet_01v8__keta_diff_25}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {2.2630378+sky130_fd_pr__pfet_01v8__ags_diff_25}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_25}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_25}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19745917+sky130_fd_pr__pfet_01v8__voff_diff_25+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_25+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_25}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.42121655+sky130_fd_pr__pfet_01v8__eta0_diff_25}
+ etab = -0.0014146465
+ dsub = 0.42114336
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.69181881+sky130_fd_pr__pfet_01v8__pclm_diff_25}
+ pdiblc1 = 0.36806399
+ pdiblc2 = 0.0066053256
+ pdiblcb = -0.025
+ drout = 0.74812414
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.3725902e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.5108411e-9
+ alpha1 = 0.0
+ beta0 = 15.614632
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_25}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_25}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_25}
+ bgidl = {1.7649271e009+sky130_fd_pr__pfet_01v8__bgidl_diff_25}
+ cgidl = {39.040404+sky130_fd_pr__pfet_01v8__cgidl_diff_25}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.568+sky130_fd_pr__pfet_01v8__kt1_diff_25}
+ kt2 = -0.1183
+ at = 60000.0
+ ute = -0.3
+ ua1 = 1.6828e-10
+ ub1 = 4.0841e-19
+ uc1 = 1.5093e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.99431+sky130_fd_pr__pfet_01v8__vth0_diff_26+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.48147074
+ k2 = {0.021329669+sky130_fd_pr__pfet_01v8__k2_diff_26}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {73792+sky130_fd_pr__pfet_01v8__vsat_diff_26}
+ ua = {-1.3677772e-009+sky130_fd_pr__pfet_01v8__ua_diff_26}
+ ub = {1.1009815e-018+sky130_fd_pr__pfet_01v8__ub_diff_26}
+ uc = -1.1898446e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_26}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0055557+sky130_fd_pr__pfet_01v8__u0_diff_26}
+ a0 = {0.90232+sky130_fd_pr__pfet_01v8__a0_diff_26}
+ keta = {-0.013964031+sky130_fd_pr__pfet_01v8__keta_diff_26}
+ a1 = 0.0
+ a2 = 0.80253166
+ ags = {0.88641503+sky130_fd_pr__pfet_01v8__ags_diff_26}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_26}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_26}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19696621+sky130_fd_pr__pfet_01v8__voff_diff_26+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4818794+sky130_fd_pr__pfet_01v8__nfactor_diff_26+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_26}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_26}
+ etab = -3.125e-5
+ dsub = 0.29198037
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62385888+sky130_fd_pr__pfet_01v8__pclm_diff_26}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.4138212
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_26}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_26}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_26}
+ bgidl = {1.2193856e009+sky130_fd_pr__pfet_01v8__bgidl_diff_26}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_26}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.50846+sky130_fd_pr__pfet_01v8__kt1_diff_26}
+ kt2 = -0.055188
+ at = 70880.0
+ ute = -0.31763
+ ua1 = 4.4497e-10
+ ub1 = 4.4717e-19
+ uc1 = 2.432e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.27 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0303+sky130_fd_pr__pfet_01v8__vth0_diff_27+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.5179279
+ k2 = {-0.00290632+sky130_fd_pr__pfet_01v8__k2_diff_27}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {71250+sky130_fd_pr__pfet_01v8__vsat_diff_27}
+ ua = {-9.8434765e-010+sky130_fd_pr__pfet_01v8__ua_diff_27}
+ ub = {8.9208454e-019+sky130_fd_pr__pfet_01v8__ub_diff_27}
+ uc = -3.5594025e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_27}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0073808+sky130_fd_pr__pfet_01v8__u0_diff_27}
+ a0 = {1.0848+sky130_fd_pr__pfet_01v8__a0_diff_27}
+ keta = {-0.0263051+sky130_fd_pr__pfet_01v8__keta_diff_27}
+ a1 = 0.0
+ a2 = 0.9
+ ags = {0.53216408+sky130_fd_pr__pfet_01v8__ags_diff_27}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_27}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_27}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20136795+sky130_fd_pr__pfet_01v8__voff_diff_27+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.7417864+sky130_fd_pr__pfet_01v8__nfactor_diff_27+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_27}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_27}
+ etab = -7.4381556
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.61751639+sky130_fd_pr__pfet_01v8__pclm_diff_27}
+ pdiblc1 = 0.37190449
+ pdiblc2 = 0.00043
+ pdiblcb = -0.00074465016
+ drout = 0.71558706
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.9355217e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.4647337e-5
+ alpha1 = 0.0
+ beta0 = 29.894997
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_27}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_27}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_27}
+ bgidl = {1.3576698e009+sky130_fd_pr__pfet_01v8__bgidl_diff_27}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_27}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.47210483+sky130_fd_pr__pfet_01v8__kt1_diff_27}
+ kt2 = -0.047360635
+ at = 90827.44
+ ute = -0.30354133
+ ua1 = 1.8739274e-9
+ ub1 = -1.1997499e-18
+ uc1 = -1.1501394e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.28 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.051+sky130_fd_pr__pfet_01v8__vth0_diff_28+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43736265
+ k2 = {0.031706452+sky130_fd_pr__pfet_01v8__k2_diff_28}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {53437.5+sky130_fd_pr__pfet_01v8__vsat_diff_28}
+ ua = {-8.6616359e-010+sky130_fd_pr__pfet_01v8__ua_diff_28}
+ ub = {8.248837e-019+sky130_fd_pr__pfet_01v8__ub_diff_28}
+ uc = -3.923953e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_28}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0077721+sky130_fd_pr__pfet_01v8__u0_diff_28}
+ a0 = {1.1863+sky130_fd_pr__pfet_01v8__a0_diff_28}
+ keta = {-0.016628379+sky130_fd_pr__pfet_01v8__keta_diff_28}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.44134013+sky130_fd_pr__pfet_01v8__ags_diff_28}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_28}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_28}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19693365+sky130_fd_pr__pfet_01v8__voff_diff_28+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4642147+sky130_fd_pr__pfet_01v8__nfactor_diff_28+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_28}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.0005+sky130_fd_pr__pfet_01v8__eta0_diff_28}
+ etab = -0.00050000043
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.40306146+sky130_fd_pr__pfet_01v8__pclm_diff_28}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00033301928
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.9955987e+8
+ pscbe2 = 8.9405959e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.152593
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_28}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_28}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_28}
+ bgidl = {1.0816056e009+sky130_fd_pr__pfet_01v8__bgidl_diff_28}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_28}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.46426465+sky130_fd_pr__pfet_01v8__kt1_diff_28}
+ kt2 = -0.043903272
+ at = 80980.356
+ ute = -0.23506459
+ ua1 = 1.6480828e-9
+ ub1 = -6.125719e-19
+ uc1 = -1.6484291e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.29 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0568+sky130_fd_pr__pfet_01v8__vth0_diff_29+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4308629
+ k2 = {0.033407718+sky130_fd_pr__pfet_01v8__k2_diff_29}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {53437.5+sky130_fd_pr__pfet_01v8__vsat_diff_29}
+ ua = {-5.5086494e-010+sky130_fd_pr__pfet_01v8__ua_diff_29}
+ ub = {5.7205917e-019+sky130_fd_pr__pfet_01v8__ub_diff_29}
+ uc = -5.9920912e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_29}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0087771+sky130_fd_pr__pfet_01v8__u0_diff_29}
+ a0 = {1.1646+sky130_fd_pr__pfet_01v8__a0_diff_29}
+ keta = {-0.011085355+sky130_fd_pr__pfet_01v8__keta_diff_29}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.28218484+sky130_fd_pr__pfet_01v8__ags_diff_29}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_29}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_29}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20189174+sky130_fd_pr__pfet_01v8__voff_diff_29+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4302911+sky130_fd_pr__pfet_01v8__nfactor_diff_29+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_29}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_29}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.43362287+sky130_fd_pr__pfet_01v8__pclm_diff_29}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00015694727
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 8.6157876e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.0385864
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_29}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_29}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.1562359e-010+sky130_fd_pr__pfet_01v8__agidl_diff_29}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_29}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_29}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.46530874+sky130_fd_pr__pfet_01v8__kt1_diff_29}
+ kt2 = -0.024824291
+ at = 093918.77
+ ute = -0.20559356
+ ua1 = 1.9942443e-9
+ ub1 = -8.2058672e-19
+ uc1 = -1.2871612e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.30 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0593+sky130_fd_pr__pfet_01v8__vth0_diff_30+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43448553
+ k2 = {0.032987346+sky130_fd_pr__pfet_01v8__k2_diff_30}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {160312.5+sky130_fd_pr__pfet_01v8__vsat_diff_30}
+ ua = {-5.6075701e-010+sky130_fd_pr__pfet_01v8__ua_diff_30}
+ ub = {5.3841446e-019+sky130_fd_pr__pfet_01v8__ub_diff_30}
+ uc = -6.6549964e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_30}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0084399+sky130_fd_pr__pfet_01v8__u0_diff_30}
+ a0 = {1.22+sky130_fd_pr__pfet_01v8__a0_diff_30}
+ keta = {0.0051290095+sky130_fd_pr__pfet_01v8__keta_diff_30}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {0.2403728+sky130_fd_pr__pfet_01v8__ags_diff_30}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_30}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_30}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613645+sky130_fd_pr__pfet_01v8__voff_diff_30+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2442058+sky130_fd_pr__pfet_01v8__nfactor_diff_30+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_30}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_30}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.0015228006+sky130_fd_pr__pfet_01v8__pclm_diff_30}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029632464
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3760948e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.6464006
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_30}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_30}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_30}
+ bgidl = {1.181082e009+sky130_fd_pr__pfet_01v8__bgidl_diff_30}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_30}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.4485+sky130_fd_pr__pfet_01v8__kt1_diff_30}
+ kt2 = -0.0075706
+ at = 90900.0
+ ute = -0.33954
+ ua1 = 1.6104e-9
+ ub1 = -5.609e-19
+ uc1 = -1.0858e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.31 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0252+sky130_fd_pr__pfet_01v8__vth0_diff_31+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.2883544
+ k2 = {-0.27784927+sky130_fd_pr__pfet_01v8__k2_diff_31}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {62851+sky130_fd_pr__pfet_01v8__vsat_diff_31}
+ ua = {-2.5066e-009+sky130_fd_pr__pfet_01v8__ua_diff_31}
+ ub = {2.147361e-018+sky130_fd_pr__pfet_01v8__ub_diff_31}
+ uc = 1.3106218e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_31}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.002831+sky130_fd_pr__pfet_01v8__u0_diff_31}
+ a0 = {0.80836322+sky130_fd_pr__pfet_01v8__a0_diff_31}
+ keta = {-0.0091058086+sky130_fd_pr__pfet_01v8__keta_diff_31}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_31}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_31}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_31}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26404672+sky130_fd_pr__pfet_01v8__voff_diff_31+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_31+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_31}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.33576108+sky130_fd_pr__pfet_01v8__eta0_diff_31}
+ etab = -0.017513367
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.32626323+sky130_fd_pr__pfet_01v8__pclm_diff_31}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -0.0030839198
+ drout = 1.0
+ pscbe1 = 7.8591361e+8
+ pscbe2 = 9.0056008e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.3771172
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_31}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_31}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_31}
+ bgidl = {1.0458447e009+sky130_fd_pr__pfet_01v8__bgidl_diff_31}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_31}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.69+sky130_fd_pr__pfet_01v8__kt1_diff_31}
+ kt2 = -0.12196
+ at = 38000.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.32 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.01+sky130_fd_pr__pfet_01v8__vth0_diff_32+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.022193
+ k2 = {-0.16868193+sky130_fd_pr__pfet_01v8__k2_diff_32}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {81122+sky130_fd_pr__pfet_01v8__vsat_diff_32}
+ ua = {-2.2782268e-009+sky130_fd_pr__pfet_01v8__ua_diff_32}
+ ub = {1.8767816e-018+sky130_fd_pr__pfet_01v8__ub_diff_32}
+ uc = 1.5507992e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_32}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0032238+sky130_fd_pr__pfet_01v8__u0_diff_32}
+ a0 = {0.53153+sky130_fd_pr__pfet_01v8__a0_diff_32}
+ keta = {-0.023377184+sky130_fd_pr__pfet_01v8__keta_diff_32}
+ a1 = 0.0
+ a2 = 0.77170379
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_32}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_32}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_32}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28237614+sky130_fd_pr__pfet_01v8__voff_diff_32+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_32+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_32}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.17082235+sky130_fd_pr__pfet_01v8__eta0_diff_32}
+ etab = -0.057223807
+ dsub = 0.28302094
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.6363737+sky130_fd_pr__pfet_01v8__pclm_diff_32}
+ pdiblc1 = 0.18660527
+ pdiblc2 = 0.0041736876
+ pdiblcb = -0.075
+ drout = 0.94973228
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.2007436e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.6052692
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_32}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_32}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.1300561e-010+sky130_fd_pr__pfet_01v8__agidl_diff_32}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_32}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_32}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5589+sky130_fd_pr__pfet_01v8__kt1_diff_32}
+ kt2 = -0.12196
+ at = 38000.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.33 pmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.96878+sky130_fd_pr__pfet_01v8__vth0_diff_33+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 0.8245821
+ k2 = {-0.098613372+sky130_fd_pr__pfet_01v8__k2_diff_33}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {88813+sky130_fd_pr__pfet_01v8__vsat_diff_33}
+ ua = {-2.0616338e-009+sky130_fd_pr__pfet_01v8__ua_diff_33}
+ ub = {1.6412578e-018+sky130_fd_pr__pfet_01v8__ub_diff_33}
+ uc = 9.6322162e-14
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_33}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0037019+sky130_fd_pr__pfet_01v8__u0_diff_33}
+ a0 = {0.65541293+sky130_fd_pr__pfet_01v8__a0_diff_33}
+ keta = {-0.081944671+sky130_fd_pr__pfet_01v8__keta_diff_33}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {2.0484732+sky130_fd_pr__pfet_01v8__ags_diff_33}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_33}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_33}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22198655+sky130_fd_pr__pfet_01v8__voff_diff_33+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_33+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_33}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.0016778392+sky130_fd_pr__pfet_01v8__eta0_diff_33}
+ etab = -0.0050335176
+ dsub = 0.41660971
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.77261114+sky130_fd_pr__pfet_01v8__pclm_diff_33}
+ pdiblc1 = 0.4223083
+ pdiblc2 = 0.010090968
+ pdiblcb = -0.075
+ drout = 0.46881029
+ pscbe1 = 7.9999646e+8
+ pscbe2 = 8.8814871e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.1381325e-9
+ alpha1 = 0.0
+ beta0 = 15.592098
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_33}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_33}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_33}
+ bgidl = {1.5623771e009+sky130_fd_pr__pfet_01v8__bgidl_diff_33}
+ cgidl = {65.986158+sky130_fd_pr__pfet_01v8__cgidl_diff_33}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5589+sky130_fd_pr__pfet_01v8__kt1_diff_33}
+ kt2 = -0.12196
+ at = 87000.0
+ ute = -0.363
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.34 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1+sky130_fd_pr__pfet_01v8__vth0_diff_34+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47538552
+ k2 = {0.024803058+sky130_fd_pr__pfet_01v8__k2_diff_34}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {79146+sky130_fd_pr__pfet_01v8__vsat_diff_34}
+ ua = {-1.3390431e-009+sky130_fd_pr__pfet_01v8__ua_diff_34}
+ ub = {1.0685272e-018+sky130_fd_pr__pfet_01v8__ub_diff_34}
+ uc = -1.3104387e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_34}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0056754+sky130_fd_pr__pfet_01v8__u0_diff_34}
+ a0 = {0.91+sky130_fd_pr__pfet_01v8__a0_diff_34}
+ keta = {-0.010198825+sky130_fd_pr__pfet_01v8__keta_diff_34}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.83892699+sky130_fd_pr__pfet_01v8__ags_diff_34}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_34}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_34}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17876326+sky130_fd_pr__pfet_01v8__voff_diff_34+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4087522+sky130_fd_pr__pfet_01v8__nfactor_diff_34+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_34}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_34}
+ etab = -6.25e-5
+ dsub = 0.29934761
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62310492+sky130_fd_pr__pfet_01v8__pclm_diff_34}
+ pdiblc1 = 0.038852787
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.1460596e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.4042378
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_34}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_34}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_34}
+ bgidl = {1.0162377e009+sky130_fd_pr__pfet_01v8__bgidl_diff_34}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_34}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.50846+sky130_fd_pr__pfet_01v8__kt1_diff_34}
+ kt2 = -0.055188
+ at = 75000.0
+ ute = -0.37025
+ ua1 = 4.5497e-10
+ ub1 = 4.1298e-19
+ uc1 = 2.432e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.35 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0185+sky130_fd_pr__pfet_01v8__vth0_diff_35+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44520413
+ k2 = {0.018979745+sky130_fd_pr__pfet_01v8__k2_diff_35}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {49081.596+sky130_fd_pr__pfet_01v8__vsat_diff_35}
+ ua = {-1.1983058e-009+sky130_fd_pr__pfet_01v8__ua_diff_35}
+ ub = {9.052489e-019+sky130_fd_pr__pfet_01v8__ub_diff_35}
+ uc = -4.4501293e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_35}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00604+sky130_fd_pr__pfet_01v8__u0_diff_35}
+ a0 = {0.92753+sky130_fd_pr__pfet_01v8__a0_diff_35}
+ keta = {-0.0079183498+sky130_fd_pr__pfet_01v8__keta_diff_35}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.63548316+sky130_fd_pr__pfet_01v8__ags_diff_35}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_35}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_35}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20198983+sky130_fd_pr__pfet_01v8__voff_diff_35+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4224191+sky130_fd_pr__pfet_01v8__nfactor_diff_35+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_35}
+ cit = 5.0e-6
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_35}
+ etab = -0.2475
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63184034+sky130_fd_pr__pfet_01v8__pclm_diff_35}
+ pdiblc1 = 0.38661844
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 0.74151816
+ pscbe1 = 7.7639675e+8
+ pscbe2 = 9.0467233e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.3542943
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_35}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_35}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.4624786e-009+sky130_fd_pr__pfet_01v8__agidl_diff_35}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_35}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_35}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.49027517+sky130_fd_pr__pfet_01v8__kt1_diff_35}
+ kt2 = -0.0628081
+ at = 59868.851
+ ute = -0.72839873
+ ua1 = -1.266648e-10
+ ub1 = 8.2317753e-19
+ uc1 = 2.7670692e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1.9995e-05 lmax = 2.0005e-05 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0212+sky130_fd_pr__pfet_01v8__vth0_diff_36+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.45790807
+ k2 = {0.018024243+sky130_fd_pr__pfet_01v8__k2_diff_36}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80156.25+sky130_fd_pr__pfet_01v8__vsat_diff_36}
+ ua = {-7.570088e-010+sky130_fd_pr__pfet_01v8__ua_diff_36}
+ ub = {5.4777974e-019+sky130_fd_pr__pfet_01v8__ub_diff_36}
+ uc = -8.5483015e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_36}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0072219031+sky130_fd_pr__pfet_01v8__u0_diff_36}
+ a0 = {1.5948701+sky130_fd_pr__pfet_01v8__a0_diff_36}
+ keta = {0.024695495+sky130_fd_pr__pfet_01v8__keta_diff_36}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {0.13602092+sky130_fd_pr__pfet_01v8__ags_diff_36}
+ b0 = {2.1073424e-024+sky130_fd_pr__pfet_01v8__b0_diff_36}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_36}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.21692555+sky130_fd_pr__pfet_01v8__voff_diff_36+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.1762342+sky130_fd_pr__pfet_01v8__nfactor_diff_36+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_36}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_36}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.00014062526+sky130_fd_pr__pfet_01v8__pclm_diff_36}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.002415402
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 6.4515428e+8
+ pscbe2 = 9.8993167e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_36}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_36}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.6391226e-010+sky130_fd_pr__pfet_01v8__agidl_diff_36}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_36}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_36}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.33852+sky130_fd_pr__pfet_01v8__kt1_diff_36}
+ kt2 = -0.058950563
+ at = 85037.625
+ ute = -0.30074
+ ua1 = 6.1946953e-10
+ ub1 = 2.4505638e-19
+ uc1 = 6.9179234e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.37 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0592+sky130_fd_pr__pfet_01v8__vth0_diff_37+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44592753
+ k2 = {0.015972271+sky130_fd_pr__pfet_01v8__k2_diff_37}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {49380.119+sky130_fd_pr__pfet_01v8__vsat_diff_37}
+ ua = {-7.2679845e-010+sky130_fd_pr__pfet_01v8__ua_diff_37}
+ ub = {5.7700106e-019+sky130_fd_pr__pfet_01v8__ub_diff_37}
+ uc = -7.5897166e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_37}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0081816+sky130_fd_pr__pfet_01v8__u0_diff_37}
+ a0 = {1.2597+sky130_fd_pr__pfet_01v8__a0_diff_37}
+ keta = {0.0022726651+sky130_fd_pr__pfet_01v8__keta_diff_37}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.36766305+sky130_fd_pr__pfet_01v8__ags_diff_37}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_37}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_37}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1989501+sky130_fd_pr__pfet_01v8__voff_diff_37+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8692119+sky130_fd_pr__pfet_01v8__nfactor_diff_37+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_37}
+ cit = 5.0e-6
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.0005+sky130_fd_pr__pfet_01v8__eta0_diff_37}
+ etab = -0.0005
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.5961172+sky130_fd_pr__pfet_01v8__pclm_diff_37}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012740962
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.4514865e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_37}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_37}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {7.0886768e-010+sky130_fd_pr__pfet_01v8__agidl_diff_37}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_37}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_37}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.4557912+sky130_fd_pr__pfet_01v8__kt1_diff_37}
+ kt2 = -0.055290049
+ at = 74171.068
+ ute = -0.81384787
+ ua1 = -2.8581502e-11
+ ub1 = 7.1990413e-19
+ uc1 = 4.3822176e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.38 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0360683+sky130_fd_pr__pfet_01v8__vth0_diff_38+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.46819224
+ k2 = {0.012171982+sky130_fd_pr__pfet_01v8__k2_diff_38}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {41389.72+sky130_fd_pr__pfet_01v8__vsat_diff_38}
+ ua = {-7.7919975e-010+sky130_fd_pr__pfet_01v8__ua_diff_38}
+ ub = {5.8244673e-019+sky130_fd_pr__pfet_01v8__ub_diff_38}
+ uc = -8.0891376e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_38}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0073118742+sky130_fd_pr__pfet_01v8__u0_diff_38}
+ a0 = {1.2673278+sky130_fd_pr__pfet_01v8__a0_diff_38}
+ keta = {0.010038944+sky130_fd_pr__pfet_01v8__keta_diff_38}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.22521628+sky130_fd_pr__pfet_01v8__ags_diff_38}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_38}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_38}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.208872+sky130_fd_pr__pfet_01v8__voff_diff_38+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8416979+sky130_fd_pr__pfet_01v8__nfactor_diff_38+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_38}
+ cit = 5.0e-6
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_38}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.61293861+sky130_fd_pr__pfet_01v8__pclm_diff_38}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00049863771
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 7.8753982e+8
+ pscbe2 = 9.4859328e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.8256686
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_38}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_38}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {8.4439949e-010+sky130_fd_pr__pfet_01v8__agidl_diff_38}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_38}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_38}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.4057912+sky130_fd_pr__pfet_01v8__kt1_diff_38}
+ kt2 = -0.055290049
+ at = 63787.0
+ ute = -0.65108
+ ua1 = -2.8581502e-11
+ ub1 = 7.1990413e-19
+ uc1 = 4.3822176e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.39 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0360683+sky130_fd_pr__pfet_01v8__vth0_diff_39+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.46819224
+ k2 = {0.012171982+sky130_fd_pr__pfet_01v8__k2_diff_39}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {41389.72+sky130_fd_pr__pfet_01v8__vsat_diff_39}
+ ua = {-7.7919975e-010+sky130_fd_pr__pfet_01v8__ua_diff_39}
+ ub = {5.8244673e-019+sky130_fd_pr__pfet_01v8__ub_diff_39}
+ uc = -8.0891376e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_39}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0073118742+sky130_fd_pr__pfet_01v8__u0_diff_39}
+ a0 = {1.2673278+sky130_fd_pr__pfet_01v8__a0_diff_39}
+ keta = {0.010038944+sky130_fd_pr__pfet_01v8__keta_diff_39}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.22521628+sky130_fd_pr__pfet_01v8__ags_diff_39}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_39}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_39}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.208872+sky130_fd_pr__pfet_01v8__voff_diff_39+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8416979+sky130_fd_pr__pfet_01v8__nfactor_diff_39+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_39}
+ cit = 5.0e-6
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_39}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.61293861+sky130_fd_pr__pfet_01v8__pclm_diff_39}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00049863771
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 7.8753982e+8
+ pscbe2 = 9.4859328e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.8256686
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_39}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_39}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {8.4439949e-010+sky130_fd_pr__pfet_01v8__agidl_diff_39}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_39}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_39}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.38852+sky130_fd_pr__pfet_01v8__kt1_diff_39}
+ kt2 = -0.058950563
+ at = 85037.625
+ ute = -0.30074
+ ua1 = 6.1946953e-10
+ ub1 = 2.4505638e-19
+ uc1 = 6.2379234e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.40 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0323+sky130_fd_pr__pfet_01v8__vth0_diff_40+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.0277986
+ k2 = {-0.19795455+sky130_fd_pr__pfet_01v8__k2_diff_40}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {105140+sky130_fd_pr__pfet_01v8__vsat_diff_40}
+ ua = {-2.4561e-009+sky130_fd_pr__pfet_01v8__ua_diff_40}
+ ub = {2.1606909e-018+sky130_fd_pr__pfet_01v8__ub_diff_40}
+ uc = 2.2568886e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_40}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0025008+sky130_fd_pr__pfet_01v8__u0_diff_40}
+ a0 = {0.87084038+sky130_fd_pr__pfet_01v8__a0_diff_40}
+ keta = {0.012330587+sky130_fd_pr__pfet_01v8__keta_diff_40}
+ a1 = 0.0
+ a2 = 0.54238276
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_40}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_40}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_40}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2787342+sky130_fd_pr__pfet_01v8__voff_diff_40+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_40+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_40}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.076984736+sky130_fd_pr__pfet_01v8__eta0_diff_40}
+ etab = -0.046584917
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.78749614+sky130_fd_pr__pfet_01v8__pclm_diff_40}
+ pdiblc1 = 0.3180521
+ pdiblc2 = 0.006885257
+ pdiblcb = -0.00014648438
+ drout = 0.90968666
+ pscbe1 = 7.9703501e+8
+ pscbe2 = 8.0953459e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.7274723
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_40}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_40}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.871786e-009+sky130_fd_pr__pfet_01v8__agidl_diff_40}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_40}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_40}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.6226+sky130_fd_pr__pfet_01v8__kt1_diff_40}
+ kt2 = -0.12
+ at = 64315.0
+ ute = -0.16211
+ ua1 = 1.3034e-10
+ ub1 = 3.7264e-19
+ uc1 = 3.8e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.41 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0373+sky130_fd_pr__pfet_01v8__vth0_diff_41+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 0.98235464
+ k2 = {-0.17228163+sky130_fd_pr__pfet_01v8__k2_diff_41}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {99337+sky130_fd_pr__pfet_01v8__vsat_diff_41}
+ ua = {-2.431704e-009+sky130_fd_pr__pfet_01v8__ua_diff_41}
+ ub = {2.0213144e-018+sky130_fd_pr__pfet_01v8__ub_diff_41}
+ uc = 7.5355966e-14
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_41}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0023496+sky130_fd_pr__pfet_01v8__u0_diff_41}
+ a0 = {1.3007+sky130_fd_pr__pfet_01v8__a0_diff_41}
+ keta = {0.060375321+sky130_fd_pr__pfet_01v8__keta_diff_41}
+ a1 = 0.0
+ a2 = 0.66860639
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_41}
+ b0 = {2.1073424e-024+sky130_fd_pr__pfet_01v8__b0_diff_41}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_41}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17771+sky130_fd_pr__pfet_01v8__voff_diff_41+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3131559+sky130_fd_pr__pfet_01v8__nfactor_diff_41+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_41}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.12366733+sky130_fd_pr__pfet_01v8__eta0_diff_41}
+ etab = -0.09888831
+ dsub = 0.26110114
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62598571+sky130_fd_pr__pfet_01v8__pclm_diff_41}
+ pdiblc1 = 0.16915343
+ pdiblc2 = 0.0033817302
+ pdiblcb = -5.7845904e-6
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.3762147
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_41}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_41}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {4.6155213e-009+sky130_fd_pr__pfet_01v8__agidl_diff_41}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_41}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_41}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.6226+sky130_fd_pr__pfet_01v8__kt1_diff_41}
+ kt2 = -0.12
+ at = 95186.0
+ ute = -0.13211
+ ua1 = 1.6553e-10
+ ub1 = 3.7264e-19
+ uc1 = 2.432e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.42 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0005+sky130_fd_pr__pfet_01v8__vth0_diff_42+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.51176178
+ k2 = {0.00019771682+sky130_fd_pr__pfet_01v8__k2_diff_42}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {57805+sky130_fd_pr__pfet_01v8__vsat_diff_42}
+ ua = {-1.6262877e-009+sky130_fd_pr__pfet_01v8__ua_diff_42}
+ ub = {1.273094e-018+sky130_fd_pr__pfet_01v8__ub_diff_42}
+ uc = -2.2175357e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_42}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.00461+sky130_fd_pr__pfet_01v8__u0_diff_42}
+ a0 = {1.2263517+sky130_fd_pr__pfet_01v8__a0_diff_42}
+ keta = {-0.033035426+sky130_fd_pr__pfet_01v8__keta_diff_42}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {1.2400293+sky130_fd_pr__pfet_01v8__ags_diff_42}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_42}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_42}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19223969+sky130_fd_pr__pfet_01v8__voff_diff_42+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8641584+sky130_fd_pr__pfet_01v8__nfactor_diff_42+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_42}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_42}
+ etab = -3.125e-6
+ dsub = 0.33687873
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.65599457+sky130_fd_pr__pfet_01v8__pclm_diff_42}
+ pdiblc1 = 0.3510864
+ pdiblc2 = 0.0018311678
+ pdiblcb = -0.025
+ drout = 0.85848102
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.2905491e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.3029989
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_42}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_42}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {6.6338926e-010+sky130_fd_pr__pfet_01v8__agidl_diff_42}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_42}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_42}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5094+sky130_fd_pr__pfet_01v8__kt1_diff_42}
+ kt2 = -0.097524
+ at = 52861.0
+ ute = -0.14338
+ ua1 = 3.9366e-10
+ ub1 = 4.6246e-19
+ uc1 = 2.432e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.43 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97494+sky130_fd_pr__pfet_01v8__vth0_diff_43+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.48496486
+ k2 = {0.012297174+sky130_fd_pr__pfet_01v8__k2_diff_43}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {66390.655+sky130_fd_pr__pfet_01v8__vsat_diff_43}
+ ua = {-1.6434761e-009+sky130_fd_pr__pfet_01v8__ua_diff_43}
+ ub = {1.2427297e-018+sky130_fd_pr__pfet_01v8__ub_diff_43}
+ uc = -2.5044847e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_43}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0042844+sky130_fd_pr__pfet_01v8__u0_diff_43}
+ a0 = {1.2214+sky130_fd_pr__pfet_01v8__a0_diff_43}
+ keta = {0.00059380239+sky130_fd_pr__pfet_01v8__keta_diff_43}
+ a1 = 0.0
+ a2 = 0.4
+ ags = {0.45174705+sky130_fd_pr__pfet_01v8__ags_diff_43}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_43}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_43}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18325928+sky130_fd_pr__pfet_01v8__voff_diff_43+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4450451+sky130_fd_pr__pfet_01v8__nfactor_diff_43+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_43}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_43}
+ etab = -0.165
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.67810107+sky130_fd_pr__pfet_01v8__pclm_diff_43}
+ pdiblc1 = 0.39050845
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 0.88837014
+ pscbe1 = 7.9879629e+8
+ pscbe2 = 9.0075561e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.9245513
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_43}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_43}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {6.2998882e-010+sky130_fd_pr__pfet_01v8__agidl_diff_43}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_43}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_43}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.51864308+sky130_fd_pr__pfet_01v8__kt1_diff_43}
+ kt2 = -0.059720037
+ at = 72802.763
+ ute = -0.180356099
+ ua1 = 1.0032102e-9
+ ub1 = -4.8656886e-19
+ uc1 = -2.5962119e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.045+sky130_fd_pr__pfet_01v8__vth0_diff_44+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44943216
+ k2 = {0.017004345+sky130_fd_pr__pfet_01v8__k2_diff_44}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {32292.293+sky130_fd_pr__pfet_01v8__vsat_diff_44}
+ ua = {-6.299923e-010+sky130_fd_pr__pfet_01v8__ua_diff_44}
+ ub = {5.6568626e-019+sky130_fd_pr__pfet_01v8__ub_diff_44}
+ uc = -6.6419472e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_44}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0083201+sky130_fd_pr__pfet_01v8__u0_diff_44}
+ a0 = {1.1618+sky130_fd_pr__pfet_01v8__a0_diff_44}
+ keta = {-0.0053050146+sky130_fd_pr__pfet_01v8__keta_diff_44}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.57074104+sky130_fd_pr__pfet_01v8__ags_diff_44}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_44}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_44}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.18907881+sky130_fd_pr__pfet_01v8__voff_diff_44+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_44+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_44}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.0005+sky130_fd_pr__pfet_01v8__eta0_diff_44}
+ etab = -0.0005
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.3006686+sky130_fd_pr__pfet_01v8__pclm_diff_44}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028889885
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.5282005e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.7149557e-12
+ alpha1 = -5.0822792e-16
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_44}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_44}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.5195639e-010+sky130_fd_pr__pfet_01v8__agidl_diff_44}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_44}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_44}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.49074474+sky130_fd_pr__pfet_01v8__kt1_diff_44}
+ kt2 = -0.057500469
+ at = 39933.378
+ ute = -0.96542388
+ ua1 = -8.8723806e-12
+ ub1 = 5.1623676e-19
+ uc1 = 4.6133748e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.45 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0123+sky130_fd_pr__pfet_01v8__vth0_diff_45+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4623874
+ k2 = {0.013868507+sky130_fd_pr__pfet_01v8__k2_diff_45}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {35932+sky130_fd_pr__pfet_01v8__vsat_diff_45}
+ ua = {-8.4255435e-010+sky130_fd_pr__pfet_01v8__ua_diff_45}
+ ub = {6.1445639e-019+sky130_fd_pr__pfet_01v8__ub_diff_45}
+ uc = -7.2682265e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_45}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0068803+sky130_fd_pr__pfet_01v8__u0_diff_45}
+ a0 = {1.2479612+sky130_fd_pr__pfet_01v8__a0_diff_45}
+ keta = {0.010639281+sky130_fd_pr__pfet_01v8__keta_diff_45}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.23404099+sky130_fd_pr__pfet_01v8__ags_diff_45}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_45}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_45}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19251341+sky130_fd_pr__pfet_01v8__voff_diff_45+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_45+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_45}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_45}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.39982968+sky130_fd_pr__pfet_01v8__pclm_diff_45}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.5793364e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.1282262e-11
+ alpha1 = 3.3623512e-17
+ beta0 = 23.665851
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_45}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_45}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_45}
+ bgidl = {1.3216319e009+sky130_fd_pr__pfet_01v8__bgidl_diff_45}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_45}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.39295+sky130_fd_pr__pfet_01v8__kt1_diff_45}
+ kt2 = -0.058527666
+ at = 62801.013
+ ute = -0.36385
+ ua1 = 3.7471e-10
+ ub1 = 4.2332524e-19
+ uc1 = -4.4399073e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.46 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0208339+sky130_fd_pr__pfet_01v8__vth0_diff_46+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47866595
+ k2 = {0.0092229355+sky130_fd_pr__pfet_01v8__k2_diff_46}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {24491.02+sky130_fd_pr__pfet_01v8__vsat_diff_46}
+ ua = {-9.0665469e-010+sky130_fd_pr__pfet_01v8__ua_diff_46}
+ ub = {7.0617665e-019+sky130_fd_pr__pfet_01v8__ub_diff_46}
+ uc = -6.8009552e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_46}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0068063633+sky130_fd_pr__pfet_01v8__u0_diff_46}
+ a0 = {1.2509318+sky130_fd_pr__pfet_01v8__a0_diff_46}
+ keta = {0.0074076058+sky130_fd_pr__pfet_01v8__keta_diff_46}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.23496304+sky130_fd_pr__pfet_01v8__ags_diff_46}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_46}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_46}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20562646+sky130_fd_pr__pfet_01v8__voff_diff_46+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4717257+sky130_fd_pr__pfet_01v8__nfactor_diff_46+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_46}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_01v8__eta0_diff_46}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.0017402344+sky130_fd_pr__pfet_01v8__pclm_diff_46}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00083787503
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 7.9009731e+8
+ pscbe2 = 9.5178184e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_46}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_46}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.1731672e-009+sky130_fd_pr__pfet_01v8__agidl_diff_46}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_46}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_46}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.52561+sky130_fd_pr__pfet_01v8__kt1_diff_46}
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.47 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0464+sky130_fd_pr__pfet_01v8__vth0_diff_47+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.2239066
+ k2 = {-0.25634724+sky130_fd_pr__pfet_01v8__k2_diff_47}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {73617+sky130_fd_pr__pfet_01v8__vsat_diff_47}
+ ua = {-2.5089e-009+sky130_fd_pr__pfet_01v8__ua_diff_47}
+ ub = {2.1633632e-018+sky130_fd_pr__pfet_01v8__ub_diff_47}
+ uc = 1.5794889e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_47}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0023446+sky130_fd_pr__pfet_01v8__u0_diff_47}
+ a0 = {0.64554208+sky130_fd_pr__pfet_01v8__a0_diff_47}
+ keta = {-0.024993345+sky130_fd_pr__pfet_01v8__keta_diff_47}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {1.875+sky130_fd_pr__pfet_01v8__ags_diff_47}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_47}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_47}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22713313+sky130_fd_pr__pfet_01v8__voff_diff_47+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_47+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_47}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.1796407+sky130_fd_pr__pfet_01v8__eta0_diff_47}
+ etab = -0.022306371
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.61751648+sky130_fd_pr__pfet_01v8__pclm_diff_47}
+ pdiblc1 = 0.1778911
+ pdiblc2 = 0.003634482
+ pdiblcb = -0.075
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.401824e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.7602198
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_47}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_47}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.5135415e-009+sky130_fd_pr__pfet_01v8__agidl_diff_47}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_47}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_47}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.64237+sky130_fd_pr__pfet_01v8__kt1_diff_47}
+ kt2 = -0.12
+ at = 58655.0
+ ute = 0.0
+ ua1 = 1.5119e-10
+ ub1 = 3.7264e-19
+ uc1 = 2.4624e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.48 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.98946+sky130_fd_pr__pfet_01v8__vth0_diff_48+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53667589
+ k2 = {0.0045054957+sky130_fd_pr__pfet_01v8__k2_diff_48}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {69720+sky130_fd_pr__pfet_01v8__vsat_diff_48}
+ ua = {-1.7951102e-009+sky130_fd_pr__pfet_01v8__ua_diff_48}
+ ub = {1.3759094e-018+sky130_fd_pr__pfet_01v8__ub_diff_48}
+ uc = -1.3087782e-11
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_48}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0038066+sky130_fd_pr__pfet_01v8__u0_diff_48}
+ a0 = {1.1042+sky130_fd_pr__pfet_01v8__a0_diff_48}
+ keta = {-0.0091972121+sky130_fd_pr__pfet_01v8__keta_diff_48}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {0.83350667+sky130_fd_pr__pfet_01v8__ags_diff_48}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_48}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_48}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17300391+sky130_fd_pr__pfet_01v8__voff_diff_48+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8632931+sky130_fd_pr__pfet_01v8__nfactor_diff_48+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_48}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_01v8__eta0_diff_48}
+ etab = -6.25e-6
+ dsub = 0.29764773
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63071024+sky130_fd_pr__pfet_01v8__pclm_diff_48}
+ pdiblc1 = 0.19617314
+ pdiblc2 = 0.00093647154
+ pdiblcb = -0.225
+ drout = 0.83538665
+ pscbe1 = 8.0e+8
+ pscbe2 = 1.0e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.058962
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_48}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_48}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.2844866e-010+sky130_fd_pr__pfet_01v8__agidl_diff_48}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_48}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_48}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.5094+sky130_fd_pr__pfet_01v8__kt1_diff_48}
+ kt2 = -0.0756
+ at = 65900.0
+ ute = -0.09202
+ ua1 = 3.1243e-10
+ ub1 = 4.7698e-19
+ uc1 = 2.432e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.49 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 6.35e-07 wmax = 6.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.96845+sky130_fd_pr__pfet_01v8__vth0_diff_49+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3315493
+ k2 = {-0.29691829+sky130_fd_pr__pfet_01v8__k2_diff_49}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {62402+sky130_fd_pr__pfet_01v8__vsat_diff_49}
+ ua = {-2.5366e-009+sky130_fd_pr__pfet_01v8__ua_diff_49}
+ ub = {2.2447373e-018+sky130_fd_pr__pfet_01v8__ub_diff_49}
+ uc = 1.4357061e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_49}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0022802+sky130_fd_pr__pfet_01v8__u0_diff_49}
+ a0 = {1.0580285+sky130_fd_pr__pfet_01v8__a0_diff_49}
+ keta = {-0.00015453568+sky130_fd_pr__pfet_01v8__keta_diff_49}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_49}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_49}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_49}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.4054369+sky130_fd_pr__pfet_01v8__voff_diff_49+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_49+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_49}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.348191+sky130_fd_pr__pfet_01v8__eta0_diff_49}
+ etab = -8.4285119e-14
+ dsub = 0.26479624
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.22269768+sky130_fd_pr__pfet_01v8__pclm_diff_49}
+ pdiblc1 = 0.00975
+ pdiblc2 = 0.000215
+ pdiblcb = -0.006154844
+ drout = 1.0
+ pscbe1 = 7.9996729e+8
+ pscbe2 = 9.0350062e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.7098269
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_49}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_49}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.7235637e-009+sky130_fd_pr__pfet_01v8__agidl_diff_49}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_49}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_49}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_49}
+ kt2 = -0.12
+ at = 41805.0
+ ute = -0.18156
+ ua1 = 1.7466e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.50 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 8.35e-07 wmax = 8.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.98654+sky130_fd_pr__pfet_01v8__vth0_diff_50+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3407728
+ k2 = {-0.27543757+sky130_fd_pr__pfet_01v8__k2_diff_50}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {54410+sky130_fd_pr__pfet_01v8__vsat_diff_50}
+ ua = {-2.5866e-009+sky130_fd_pr__pfet_01v8__ua_diff_50}
+ ub = {2.1888883e-018+sky130_fd_pr__pfet_01v8__ub_diff_50}
+ uc = 1.5441351e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_50}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0019711+sky130_fd_pr__pfet_01v8__u0_diff_50}
+ a0 = {1.0472628+sky130_fd_pr__pfet_01v8__a0_diff_50}
+ keta = {0.0966341+sky130_fd_pr__pfet_01v8__keta_diff_50}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {0.57891652+sky130_fd_pr__pfet_01v8__ags_diff_50}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_50}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_50}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.32071362+sky130_fd_pr__pfet_01v8__voff_diff_50+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_50+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_50}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.40158237+sky130_fd_pr__pfet_01v8__eta0_diff_50}
+ etab = -0.041512856
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.28533384+sky130_fd_pr__pfet_01v8__pclm_diff_50}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.4414063e-5
+ drout = 1.0
+ pscbe1 = 7.690463e+8
+ pscbe2 = 8.8014656e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.2607902
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_50}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_50}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.2137475e-010+sky130_fd_pr__pfet_01v8__agidl_diff_50}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_50}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_50}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_50}
+ kt2 = -0.12
+ at = 21109.0
+ ute = -0.21243
+ ua1 = 1.0762e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.51 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.645e-06 wmax = 1.655e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.02+sky130_fd_pr__pfet_01v8__vth0_diff_51+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3255051
+ k2 = {-0.28016116+sky130_fd_pr__pfet_01v8__k2_diff_51}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {59524+sky130_fd_pr__pfet_01v8__vsat_diff_51}
+ ua = {-2.4816e-009+sky130_fd_pr__pfet_01v8__ua_diff_51}
+ ub = {2.1055982e-018+sky130_fd_pr__pfet_01v8__ub_diff_51}
+ uc = 9.1597053e-14
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_51}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0024424+sky130_fd_pr__pfet_01v8__u0_diff_51}
+ a0 = {0.80890904+sky130_fd_pr__pfet_01v8__a0_diff_51}
+ keta = {0.027840733+sky130_fd_pr__pfet_01v8__keta_diff_51}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_51}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_51}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_51}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.27372667+sky130_fd_pr__pfet_01v8__voff_diff_51+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_51+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_51}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.3010182+sky130_fd_pr__pfet_01v8__eta0_diff_51}
+ etab = -0.035338434
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.47998966+sky130_fd_pr__pfet_01v8__pclm_diff_51}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.4222865e-5
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3226724e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.537679
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_51}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_51}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.8211658e-010+sky130_fd_pr__pfet_01v8__agidl_diff_51}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_51}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_51}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_51}
+ kt2 = -0.12
+ at = 39225.0
+ ute = -0.21243
+ ua1 = 1.6473e-10
+ ub1 = 3.6891e-19
+ uc1 = 6.4484e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.52 pmos
* DC IV MOS Parameters
+ lmin = 1.65e-07 lmax = 1.75e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0323+sky130_fd_pr__pfet_01v8__vth0_diff_40+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.0277986
+ k2 = {-0.19795455+sky130_fd_pr__pfet_01v8__k2_diff_40}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {105140+sky130_fd_pr__pfet_01v8__vsat_diff_40}
+ ua = {-2.4561e-009+sky130_fd_pr__pfet_01v8__ua_diff_40}
+ ub = {2.1606909e-018+sky130_fd_pr__pfet_01v8__ub_diff_40}
+ uc = 2.2568886e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_40}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0025008+sky130_fd_pr__pfet_01v8__u0_diff_40}
+ a0 = {0.87084038+sky130_fd_pr__pfet_01v8__a0_diff_40}
+ keta = {0.012330587+sky130_fd_pr__pfet_01v8__keta_diff_40}
+ a1 = 0.0
+ a2 = 0.54238276
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_40}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_40}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_40}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2787342+sky130_fd_pr__pfet_01v8__voff_diff_40+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_40+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_40}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.076984736+sky130_fd_pr__pfet_01v8__eta0_diff_40}
+ etab = -0.046584917
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.78749614+sky130_fd_pr__pfet_01v8__pclm_diff_40}
+ pdiblc1 = 0.3180521
+ pdiblc2 = 0.006885257
+ pdiblcb = -0.00014648438
+ drout = 0.90968666
+ pscbe1 = 7.9703501e+8
+ pscbe2 = 8.0953459e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.7274723
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_40}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_40}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.871786e-009+sky130_fd_pr__pfet_01v8__agidl_diff_40}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_40}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_40}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.6226+sky130_fd_pr__pfet_01v8__kt1_diff_40}
+ kt2 = -0.12
+ at = 64315.0
+ ute = -0.16211
+ ua1 = 1.3034e-10
+ ub1 = 3.7264e-19
+ uc1 = 3.8e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.53 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0464+sky130_fd_pr__pfet_01v8__vth0_diff_47+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.2239066
+ k2 = {-0.25634724+sky130_fd_pr__pfet_01v8__k2_diff_47}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {73617+sky130_fd_pr__pfet_01v8__vsat_diff_47}
+ ua = {-2.5089e-009+sky130_fd_pr__pfet_01v8__ua_diff_47}
+ ub = {2.1633632e-018+sky130_fd_pr__pfet_01v8__ub_diff_47}
+ uc = 1.5794889e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_47}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0023446+sky130_fd_pr__pfet_01v8__u0_diff_47}
+ a0 = {0.64554208+sky130_fd_pr__pfet_01v8__a0_diff_47}
+ keta = {-0.024993345+sky130_fd_pr__pfet_01v8__keta_diff_47}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {1.875+sky130_fd_pr__pfet_01v8__ags_diff_47}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_47}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_47}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22713313+sky130_fd_pr__pfet_01v8__voff_diff_47+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_47+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_47}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.1796407+sky130_fd_pr__pfet_01v8__eta0_diff_47}
+ etab = -0.022306371
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.61751648+sky130_fd_pr__pfet_01v8__pclm_diff_47}
+ pdiblc1 = 0.1778911
+ pdiblc2 = 0.003634482
+ pdiblcb = -0.075
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.401824e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.7602198
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_47}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_47}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.5135415e-009+sky130_fd_pr__pfet_01v8__agidl_diff_47}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_47}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_47}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.64237+sky130_fd_pr__pfet_01v8__kt1_diff_47}
+ kt2 = -0.12
+ at = 58655.0
+ ute = 0.0
+ ua1 = 1.5119e-10
+ ub1 = 3.7264e-19
+ uc1 = 2.4624e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.54 pmos
* DC IV MOS Parameters
+ lmin = 1.65e-07 lmax = 1.75e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.0464+sky130_fd_pr__pfet_01v8__vth0_diff_47+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.2239066
+ k2 = {-0.25634724+sky130_fd_pr__pfet_01v8__k2_diff_47}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {73617+sky130_fd_pr__pfet_01v8__vsat_diff_47}
+ ua = {-2.5089e-009+sky130_fd_pr__pfet_01v8__ua_diff_47}
+ ub = {2.1633632e-018+sky130_fd_pr__pfet_01v8__ub_diff_47}
+ uc = 1.5794889e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_47}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0023446+sky130_fd_pr__pfet_01v8__u0_diff_47}
+ a0 = {0.64554208+sky130_fd_pr__pfet_01v8__a0_diff_47}
+ keta = {-0.024993345+sky130_fd_pr__pfet_01v8__keta_diff_47}
+ a1 = 0.0
+ a2 = 0.8
+ ags = {1.875+sky130_fd_pr__pfet_01v8__ags_diff_47}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_47}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_47}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22713313+sky130_fd_pr__pfet_01v8__voff_diff_47+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_47+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_47}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.1796407+sky130_fd_pr__pfet_01v8__eta0_diff_47}
+ etab = -0.022306371
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.61751648+sky130_fd_pr__pfet_01v8__pclm_diff_47}
+ pdiblc1 = 0.1778911
+ pdiblc2 = 0.003634482
+ pdiblcb = -0.075
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.401824e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.7602198
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_47}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_47}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.5135415e-009+sky130_fd_pr__pfet_01v8__agidl_diff_47}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_47}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_47}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.64237+sky130_fd_pr__pfet_01v8__kt1_diff_47}
+ kt2 = -0.12
+ at = 58655.0
+ ute = 0.0
+ ua1 = 1.5119e-10
+ ub1 = 3.7264e-19
+ uc1 = 2.4624e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.55 pmos
* DC IV MOS Parameters
+ lmin = 1.65e-07 lmax = 1.75e-07 wmin = 6.35e-07 wmax = 6.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.96845+sky130_fd_pr__pfet_01v8__vth0_diff_49+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3315493
+ k2 = {-0.29691829+sky130_fd_pr__pfet_01v8__k2_diff_49}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {62402+sky130_fd_pr__pfet_01v8__vsat_diff_49}
+ ua = {-2.5366e-009+sky130_fd_pr__pfet_01v8__ua_diff_49}
+ ub = {2.2447373e-018+sky130_fd_pr__pfet_01v8__ub_diff_49}
+ uc = 1.4357061e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_49}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0022802+sky130_fd_pr__pfet_01v8__u0_diff_49}
+ a0 = {1.0580285+sky130_fd_pr__pfet_01v8__a0_diff_49}
+ keta = {-0.00015453568+sky130_fd_pr__pfet_01v8__keta_diff_49}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_49}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_49}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_49}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.4054369+sky130_fd_pr__pfet_01v8__voff_diff_49+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_49+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_49}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.348191+sky130_fd_pr__pfet_01v8__eta0_diff_49}
+ etab = -8.4285119e-14
+ dsub = 0.26479624
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.22269768+sky130_fd_pr__pfet_01v8__pclm_diff_49}
+ pdiblc1 = 0.00975
+ pdiblc2 = 0.000215
+ pdiblcb = -0.006154844
+ drout = 1.0
+ pscbe1 = 7.9996729e+8
+ pscbe2 = 9.0350062e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.7098269
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_49}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_49}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.7235637e-009+sky130_fd_pr__pfet_01v8__agidl_diff_49}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_49}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_49}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_49}
+ kt2 = -0.12
+ at = 41805.0
+ ute = -0.18156
+ ua1 = 1.7466e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.56 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 6.35e-07 wmax = 6.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.96845+sky130_fd_pr__pfet_01v8__vth0_diff_49+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3315493
+ k2 = {-0.29691829+sky130_fd_pr__pfet_01v8__k2_diff_49}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {62402+sky130_fd_pr__pfet_01v8__vsat_diff_49}
+ ua = {-2.5366e-009+sky130_fd_pr__pfet_01v8__ua_diff_49}
+ ub = {2.2447373e-018+sky130_fd_pr__pfet_01v8__ub_diff_49}
+ uc = 1.4357061e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_49}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0022802+sky130_fd_pr__pfet_01v8__u0_diff_49}
+ a0 = {1.0580285+sky130_fd_pr__pfet_01v8__a0_diff_49}
+ keta = {-0.00015453568+sky130_fd_pr__pfet_01v8__keta_diff_49}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_49}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_49}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_49}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.4054369+sky130_fd_pr__pfet_01v8__voff_diff_49+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_49+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_49}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.348191+sky130_fd_pr__pfet_01v8__eta0_diff_49}
+ etab = -8.4285119e-14
+ dsub = 0.26479624
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.22269768+sky130_fd_pr__pfet_01v8__pclm_diff_49}
+ pdiblc1 = 0.00975
+ pdiblc2 = 0.000215
+ pdiblcb = -0.006154844
+ drout = 1.0
+ pscbe1 = 7.9996729e+8
+ pscbe2 = 9.0350062e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.7098269
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_49}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_49}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.7235637e-009+sky130_fd_pr__pfet_01v8__agidl_diff_49}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_49}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_49}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_49}
+ kt2 = -0.12
+ at = 41805.0
+ ute = -0.18156
+ ua1 = 1.7466e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.57 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 8.35e-07 wmax = 8.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.98654+sky130_fd_pr__pfet_01v8__vth0_diff_50+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3407728
+ k2 = {-0.27543757+sky130_fd_pr__pfet_01v8__k2_diff_50}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {54410+sky130_fd_pr__pfet_01v8__vsat_diff_50}
+ ua = {-2.5866e-009+sky130_fd_pr__pfet_01v8__ua_diff_50}
+ ub = {2.1888883e-018+sky130_fd_pr__pfet_01v8__ub_diff_50}
+ uc = 1.5441351e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_50}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0019711+sky130_fd_pr__pfet_01v8__u0_diff_50}
+ a0 = {1.0472628+sky130_fd_pr__pfet_01v8__a0_diff_50}
+ keta = {0.0966341+sky130_fd_pr__pfet_01v8__keta_diff_50}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {0.57891652+sky130_fd_pr__pfet_01v8__ags_diff_50}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_50}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_50}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.32071362+sky130_fd_pr__pfet_01v8__voff_diff_50+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_50+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_50}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.40158237+sky130_fd_pr__pfet_01v8__eta0_diff_50}
+ etab = -0.041512856
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.28533384+sky130_fd_pr__pfet_01v8__pclm_diff_50}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.4414063e-5
+ drout = 1.0
+ pscbe1 = 7.690463e+8
+ pscbe2 = 8.8014656e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.2607902
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_50}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_50}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.2137475e-010+sky130_fd_pr__pfet_01v8__agidl_diff_50}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_50}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_50}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_50}
+ kt2 = -0.12
+ at = 21109.0
+ ute = -0.21243
+ ua1 = 1.0762e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.58 pmos
* DC IV MOS Parameters
+ lmin = 1.65e-07 lmax = 1.75e-07 wmin = 8.35e-07 wmax = 8.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.98654+sky130_fd_pr__pfet_01v8__vth0_diff_50+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.3407728
+ k2 = {-0.27543757+sky130_fd_pr__pfet_01v8__k2_diff_50}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {54410+sky130_fd_pr__pfet_01v8__vsat_diff_50}
+ ua = {-2.5866e-009+sky130_fd_pr__pfet_01v8__ua_diff_50}
+ ub = {2.1888883e-018+sky130_fd_pr__pfet_01v8__ub_diff_50}
+ uc = 1.5441351e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_50}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0019711+sky130_fd_pr__pfet_01v8__u0_diff_50}
+ a0 = {1.0472628+sky130_fd_pr__pfet_01v8__a0_diff_50}
+ keta = {0.0966341+sky130_fd_pr__pfet_01v8__keta_diff_50}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {0.57891652+sky130_fd_pr__pfet_01v8__ags_diff_50}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_50}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_50}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.32071362+sky130_fd_pr__pfet_01v8__voff_diff_50+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_50+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_50}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.40158237+sky130_fd_pr__pfet_01v8__eta0_diff_50}
+ etab = -0.041512856
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.28533384+sky130_fd_pr__pfet_01v8__pclm_diff_50}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.4414063e-5
+ drout = 1.0
+ pscbe1 = 7.690463e+8
+ pscbe2 = 8.8014656e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.2607902
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_50}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_50}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.2137475e-010+sky130_fd_pr__pfet_01v8__agidl_diff_50}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_50}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_50}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_50}
+ kt2 = -0.12
+ at = 21109.0
+ ute = -0.21243
+ ua1 = 1.0762e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.59 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 1.115e-06 wmax = 1.125e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.95759+sky130_fd_pr__pfet_01v8__vth0_diff_7+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.1286524
+ k2 = {-0.20642701+sky130_fd_pr__pfet_01v8__k2_diff_7}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {81677+sky130_fd_pr__pfet_01v8__vsat_diff_7}
+ ua = {-2.3466042e-009+sky130_fd_pr__pfet_01v8__ua_diff_7}
+ ub = {1.9914931e-018+sky130_fd_pr__pfet_01v8__ub_diff_7}
+ uc = 2.2913949e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_7}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0027565+sky130_fd_pr__pfet_01v8__u0_diff_7}
+ a0 = {1.087+sky130_fd_pr__pfet_01v8__a0_diff_7}
+ keta = {0.027122826+sky130_fd_pr__pfet_01v8__keta_diff_7}
+ a1 = 0.0
+ a2 = 0.68678659
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_7}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_7}
+ b1 = {2.1073424e-024+sky130_fd_pr__pfet_01v8__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.24161658+sky130_fd_pr__pfet_01v8__voff_diff_7+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_7+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_7}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.21136947+sky130_fd_pr__pfet_01v8__eta0_diff_7}
+ etab = -0.031554764
+ dsub = 0.26948731
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62205899+sky130_fd_pr__pfet_01v8__pclm_diff_7}
+ pdiblc1 = 0.15224245
+ pdiblc2 = 0.0023148811
+ pdiblcb = -0.075
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3883381e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.7923713
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_7}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_7}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_7}
+ bgidl = {1.0029534e009+sky130_fd_pr__pfet_01v8__bgidl_diff_7}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_7}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.63808+sky130_fd_pr__pfet_01v8__kt1_diff_7}
+ kt2 = -0.12
+ at = 59144.0
+ ute = -0.21616
+ ua1 = 1.505e-10
+ ub1 = 4.39e-19
+ uc1 = 9.4135e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.60 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 1.255e-06 wmax = 1.265e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.95759+sky130_fd_pr__pfet_01v8__vth0_diff_7+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.1286524
+ k2 = {-0.20642701+sky130_fd_pr__pfet_01v8__k2_diff_7}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {81677+sky130_fd_pr__pfet_01v8__vsat_diff_7}
+ ua = {-2.3466042e-009+sky130_fd_pr__pfet_01v8__ua_diff_7}
+ ub = {1.9914931e-018+sky130_fd_pr__pfet_01v8__ub_diff_7}
+ uc = 2.2913949e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_7}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0027565+sky130_fd_pr__pfet_01v8__u0_diff_7}
+ a0 = {1.087+sky130_fd_pr__pfet_01v8__a0_diff_7}
+ keta = {0.027122826+sky130_fd_pr__pfet_01v8__keta_diff_7}
+ a1 = 0.0
+ a2 = 0.68678659
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_7}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_7}
+ b1 = {2.1073424e-024+sky130_fd_pr__pfet_01v8__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.24161658+sky130_fd_pr__pfet_01v8__voff_diff_7+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.9+sky130_fd_pr__pfet_01v8__nfactor_diff_7+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_7}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.21136947+sky130_fd_pr__pfet_01v8__eta0_diff_7}
+ etab = -0.031554764
+ dsub = 0.26948731
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.62205899+sky130_fd_pr__pfet_01v8__pclm_diff_7}
+ pdiblc1 = 0.15224245
+ pdiblc2 = 0.0023148811
+ pdiblcb = -0.075
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3883381e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.7923713
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_7}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_7}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-010+sky130_fd_pr__pfet_01v8__agidl_diff_7}
+ bgidl = {1.0029534e009+sky130_fd_pr__pfet_01v8__bgidl_diff_7}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_7}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.63808+sky130_fd_pr__pfet_01v8__kt1_diff_7}
+ kt2 = -0.12
+ at = 59144.0
+ ute = -0.21616
+ ua1 = 1.505e-10
+ ub1 = 4.39e-19
+ uc1 = 9.4135e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.61 pmos
* DC IV MOS Parameters
+ lmin = 1.65e-07 lmax = 1.75e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97755+sky130_fd_pr__pfet_01v8__vth0_diff_6+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.4974388
+ k2 = {-0.34240453+sky130_fd_pr__pfet_01v8__k2_diff_6}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {55335+sky130_fd_pr__pfet_01v8__vsat_diff_6}
+ ua = {-2.5669e-009+sky130_fd_pr__pfet_01v8__ua_diff_6}
+ ub = {2.1902542e-018+sky130_fd_pr__pfet_01v8__ub_diff_6}
+ uc = 2.3206046e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_6}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0020949+sky130_fd_pr__pfet_01v8__u0_diff_6}
+ a0 = {0.72595373+sky130_fd_pr__pfet_01v8__a0_diff_6}
+ keta = {-0.0003767501+sky130_fd_pr__pfet_01v8__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_6}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_6}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28041511+sky130_fd_pr__pfet_01v8__voff_diff_6+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.892779+sky130_fd_pr__pfet_01v8__nfactor_diff_6+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_6}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.34230525+sky130_fd_pr__pfet_01v8__eta0_diff_6}
+ etab = -1.1566507e-13
+ dsub = 0.26628854
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.45374464+sky130_fd_pr__pfet_01v8__pclm_diff_6}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.4414063e-5
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3761341e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.2512308
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.1989212e-010+sky130_fd_pr__pfet_01v8__agidl_diff_6}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_6}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_6}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_6}
+ kt2 = -0.12
+ at = 21109.0
+ ute = -0.21243
+ ua1 = 1.0762e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.62 pmos
* DC IV MOS Parameters
+ lmin = 1.65e-07 lmax = 1.75e-07 wmin = 1.115e-06 wmax = 1.125e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97755+sky130_fd_pr__pfet_01v8__vth0_diff_6+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.4974388
+ k2 = {-0.34240453+sky130_fd_pr__pfet_01v8__k2_diff_6}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {55335+sky130_fd_pr__pfet_01v8__vsat_diff_6}
+ ua = {-2.5669e-009+sky130_fd_pr__pfet_01v8__ua_diff_6}
+ ub = {2.1902542e-018+sky130_fd_pr__pfet_01v8__ub_diff_6}
+ uc = 2.3206046e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_6}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0020949+sky130_fd_pr__pfet_01v8__u0_diff_6}
+ a0 = {0.72595373+sky130_fd_pr__pfet_01v8__a0_diff_6}
+ keta = {-0.0003767501+sky130_fd_pr__pfet_01v8__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_6}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_6}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28041511+sky130_fd_pr__pfet_01v8__voff_diff_6+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.892779+sky130_fd_pr__pfet_01v8__nfactor_diff_6+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_6}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.34230525+sky130_fd_pr__pfet_01v8__eta0_diff_6}
+ etab = -1.1566507e-13
+ dsub = 0.26628854
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.45374464+sky130_fd_pr__pfet_01v8__pclm_diff_6}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.4414063e-5
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3761341e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.2512308
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.1989212e-010+sky130_fd_pr__pfet_01v8__agidl_diff_6}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_6}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_6}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_6}
+ kt2 = -0.12
+ at = 21109.0
+ ute = -0.21243
+ ua1 = 1.0762e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.63 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 1.675e-06 wmax = 1.685e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.004+sky130_fd_pr__pfet_01v8__vth0_diff_16+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.0376715
+ k2 = {-0.17335648+sky130_fd_pr__pfet_01v8__k2_diff_16}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {88456+sky130_fd_pr__pfet_01v8__vsat_diff_16}
+ ua = {-2.2421727e-009+sky130_fd_pr__pfet_01v8__ua_diff_16}
+ ub = {1.8536584e-018+sky130_fd_pr__pfet_01v8__ub_diff_16}
+ uc = 2.5234343e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_16}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0029971+sky130_fd_pr__pfet_01v8__u0_diff_16}
+ a0 = {0.89088+sky130_fd_pr__pfet_01v8__a0_diff_16}
+ keta = {0.023895141+sky130_fd_pr__pfet_01v8__keta_diff_16}
+ a1 = 0.0
+ a2 = 0.67187683
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_16}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_16}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_16}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22630768+sky130_fd_pr__pfet_01v8__voff_diff_16+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.7534082+sky130_fd_pr__pfet_01v8__nfactor_diff_16+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_16}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.18201237+sky130_fd_pr__pfet_01v8__eta0_diff_16}
+ etab = -0.078353952
+ dsub = 0.27170577
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63088962+sky130_fd_pr__pfet_01v8__pclm_diff_16}
+ pdiblc1 = 0.18080115
+ pdiblc2 = 0.0040267418
+ pdiblcb = -0.0001934424
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.4769552e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.580652
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_16}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_16}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.0157032e-010+sky130_fd_pr__pfet_01v8__agidl_diff_16}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_16}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_16}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.598+sky130_fd_pr__pfet_01v8__kt1_diff_16}
+ kt2 = -0.12196
+ at = 68317.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.64 pmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 1.995e-06 wmax = 2.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1.004+sky130_fd_pr__pfet_01v8__vth0_diff_16+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.0376715
+ k2 = {-0.17335648+sky130_fd_pr__pfet_01v8__k2_diff_16}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {88456+sky130_fd_pr__pfet_01v8__vsat_diff_16}
+ ua = {-2.2421727e-009+sky130_fd_pr__pfet_01v8__ua_diff_16}
+ ub = {1.8536584e-018+sky130_fd_pr__pfet_01v8__ub_diff_16}
+ uc = 2.5234343e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_16}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0029971+sky130_fd_pr__pfet_01v8__u0_diff_16}
+ a0 = {0.89088+sky130_fd_pr__pfet_01v8__a0_diff_16}
+ keta = {0.023895141+sky130_fd_pr__pfet_01v8__keta_diff_16}
+ a1 = 0.0
+ a2 = 0.67187683
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_16}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_16}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_16}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.22630768+sky130_fd_pr__pfet_01v8__voff_diff_16+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.7534082+sky130_fd_pr__pfet_01v8__nfactor_diff_16+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_16}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.18201237+sky130_fd_pr__pfet_01v8__eta0_diff_16}
+ etab = -0.078353952
+ dsub = 0.27170577
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.63088962+sky130_fd_pr__pfet_01v8__pclm_diff_16}
+ pdiblc1 = 0.18080115
+ pdiblc2 = 0.0040267418
+ pdiblcb = -0.0001934424
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.4769552e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.580652
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_16}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_16}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.0157032e-010+sky130_fd_pr__pfet_01v8__agidl_diff_16}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_16}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_16}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.598+sky130_fd_pr__pfet_01v8__kt1_diff_16}
+ kt2 = -0.12196
+ at = 68317.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.65 pmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.115e-06 wmax = 1.125e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {-1.3994e-008+sky130_fd_pr__pfet_01v8__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {7.3039e-009+sky130_fd_pr__pfet_01v8__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.23e-009*sky130_fd_pr__pfet_01v8__toxe_mult+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.23e-09*sky130_fd_pr__pfet_01v8__toxe_mult*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_01v8__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97755+sky130_fd_pr__pfet_01v8__vth0_diff_6+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))}
+ k1 = 1.4974388
+ k2 = {-0.34240453+sky130_fd_pr__pfet_01v8__k2_diff_6}
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {55335+sky130_fd_pr__pfet_01v8__vsat_diff_6}
+ ua = {-2.5669e-009+sky130_fd_pr__pfet_01v8__ua_diff_6}
+ ub = {2.1902542e-018+sky130_fd_pr__pfet_01v8__ub_diff_6}
+ uc = 2.3206046e-13
+ rdsw = {547.88+sky130_fd_pr__pfet_01v8__rdsw_diff_6}
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = {0.0020949+sky130_fd_pr__pfet_01v8__u0_diff_6}
+ a0 = {0.72595373+sky130_fd_pr__pfet_01v8__a0_diff_6}
+ keta = {-0.0003767501+sky130_fd_pr__pfet_01v8__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.9995
+ ags = {1.25+sky130_fd_pr__pfet_01v8__ags_diff_6}
+ b0 = {0+sky130_fd_pr__pfet_01v8__b0_diff_6}
+ b1 = {0+sky130_fd_pr__pfet_01v8__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28041511+sky130_fd_pr__pfet_01v8__voff_diff_6+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))}
+ nfactor = {1.892779+sky130_fd_pr__pfet_01v8__nfactor_diff_6+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_01v8__tvoff_diff_6}
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = {0.34230525+sky130_fd_pr__pfet_01v8__eta0_diff_6}
+ etab = -1.1566507e-13
+ dsub = 0.26628854
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.45374464+sky130_fd_pr__pfet_01v8__pclm_diff_6}
+ pdiblc1 = 0.0195
+ pdiblc2 = 0.00043
+ pdiblcb = -2.4414063e-5
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 9.3761341e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.2512308
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_01v8__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_01v8__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.1989212e-010+sky130_fd_pr__pfet_01v8__agidl_diff_6}
+ bgidl = {1e009+sky130_fd_pr__pfet_01v8__bgidl_diff_6}
+ cgidl = {300+sky130_fd_pr__pfet_01v8__cgidl_diff_6}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = {-0.70976+sky130_fd_pr__pfet_01v8__kt1_diff_6}
+ kt2 = -0.12
+ at = 21109.0
+ ute = -0.21243
+ ua1 = 1.0762e-10
+ ub1 = 3.6891e-19
+ uc1 = 7.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgso = {5.5e-11*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_01v8__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {-3e-09+sky130_fd_pr__pfet_01v8__dlc_diff+sky130_fd_pr__pfet_01v8__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_01v8__dwc_diff}
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00074079*sky130_fd_pr__pfet_01v8__ajunction_mult}
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = {9.88e-011*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = {2.3894e-010*sky130_fd_pr__pfet_01v8__pjunction_mult}
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_01v8
