* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_01v8_hvt d g s b
+ 
.param  l = 1u w = 1u ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 nf = 1.0
msky130_fd_pr__pfet_01v8_hvt d g s b sky130_fd_pr__pfet_01v8_hvt__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
.model sky130_fd_pr__pfet_01v8_hvt__model.0 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.1097881+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43657182
+ k2 = 0.029080988
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.23239888+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3940676+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.014934398
+ ua = -5.7327697e-10
+ ub = 1.80325173e-18
+ uc = -7.7670696e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 200000.0
+ a0 = 1.477815
+ ags = 0.4141498
+ a1 = 0.0
+ a2 = 1.0
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.013169082
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.075489662
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0036275994
+ pdiblcb = -9.5744039e-5
+ drout = 0.56
+ pscbe1 = 746475130.0
+ pscbe2 = 9.5049925e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.7923891
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1154444600.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.44169
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.30066
+ ua1 = 2.2116e-9
+ ub1 = -7.9359e-19
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.1 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.1097881+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43657182
+ k2 = 0.029080988
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.23239888+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3940676+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.014934398
+ ua = -5.7327697e-10
+ ub = 1.80325173e-18
+ uc = -7.7670696e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 200000.0
+ a0 = 1.477815
+ ags = 0.4141498
+ a1 = 0.0
+ a2 = 1.0
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.013169082
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.075489662
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0036275994
+ pdiblcb = -9.5744039e-5
+ drout = 0.56
+ pscbe1 = 746475130.0
+ pscbe2 = 9.5049925e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.7923891
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1154444600.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.44169
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.30066
+ ua1 = 2.2116e-9
+ ub1 = -7.9359e-19
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.2 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.109098583e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.515630273e-09 wvth0 = -6.896985593e-08 pvth0 = 5.517081546e-13
+ k1 = 4.360518816e-01 lk1 = 4.159125175e-09 wk1 = 5.200752225e-08 pk1 = -4.160219524e-13
+ k2 = 2.942226684e-02 lk2 = -2.729979878e-09 wk2 = -3.413686370e-08 pk2 = 2.730698190e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.322912521e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.609437151e-10 wvoff = -1.076561717e-08 pvoff = 8.611702466e-14
+ nfactor = {1.392604281e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.170547974e-08 wnfactor = 1.463704439e-07 pnfactor = -1.170855969e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.492091026e-02 lu0 = 1.078919906e-10 wu0 = 1.349128690e-09 pu0 = -1.079203791e-14
+ ua = -5.709003964e-10 lua = -1.901084234e-17 wua = -2.377198964e-16 pua = 1.901584447e-21
+ ub = 1.796796757e-18 lub = 5.163503919e-26 wub = 6.456671382e-25 pub = -5.164862540e-30
+ uc = -7.712280941e-11 luc = -4.382690050e-18 wuc = -5.480307532e-17 puc = 4.383843223e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.943888537e+05 lvsat = 4.488504638e-02 wvsat = 5.612622726e-01 pvsat = -4.489685653e-6
+ a0 = 1.500781002e+00 la0 = -1.837111358e-07 wa0 = -2.297204479e-06 pa0 = 1.837594739e-11
+ ags = 4.342779995e-01 lags = -1.610108014e-07 wags = -2.013349559e-06 pags = 1.610531666e-11
+ a1 = 0.0
+ a2 = 9.848831835e-01 la2 = 1.208434283e-07 wa2 = 1.511079139e-06 pa2 = -1.208752247e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.635766497e-02 lketa = 2.550632012e-08 wketa = 3.189421946e-07 pketa = -2.551303134e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.175886361e-01 lpclm = -3.367608502e-07 wpclm = -4.211005121e-06 ppclm = 3.368494588e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.389690386e-03 lpdiblc2 = 1.903097248e-09 wpdiblc2 = 2.379716125e-08 ppdiblc2 = -1.903597991e-13
+ pdiblcb = -1.467572422e-04 lpdiblcb = 4.080681306e-10 wpdiblcb = 5.102662576e-09 ppdiblcb = -4.081755015e-14
+ drout = 0.56
+ pscbe1 = 7.505182841e+08 lpscbe1 = -3.234226108e+01 wpscbe1 = -4.044217934e+02 ppscbe1 = 3.235077097e-3
+ pscbe2 = 9.463114205e-09 lpscbe2 = 3.349955791e-16 wpscbe2 = 4.188931397e-15 ppscbe2 = -3.350837231e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.831973673e+00 lbeta0 = -3.166474873e-07 wbeta0 = -3.959498824e-06 pbeta0 = 3.167308036e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.034247778e-10 lagidl = -2.739570492e-17 wagidl = -3.425678894e-16 pagidl = 2.740291328e-21
+ bgidl = 1.142778186e+09 lbgidl = 9.332274090e+01 wbgidl = 1.166948413e+03 pbgidl = -9.334729598e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.425035427e-01 lkt1 = 6.507744004e-09 wkt1 = 8.137568041e-08 pkt1 = -6.509456321e-13
+ kt2 = -3.814115779e-02 lkt2 = 1.441129940e-09 wkt2 = 1.802051976e-08 pkt2 = -1.441509130e-13
+ at = 1.982944345e+04 lat = -1.586209729e-01 wat = -1.983466097e+00 pat = 1.586627093e-5
+ ute = -3.004779538e-01 lute = -1.456236123e-09 wute = -1.820941409e-08 pute = 1.456619288e-13
+ ua1 = 2.227221229e-09 lua1 = -1.249583528e-16 wua1 = -1.562533956e-15 pua1 = 1.249912319e-20
+ ub1 = -8.067509612e-19 lub1 = 1.052780165e-25 wub1 = 1.316442414e-24 pub1 = -1.053057173e-29
+ uc1 = 1.211394313e-10 luc1 = -1.031450233e-17 wuc1 = -1.289770533e-16 puc1 = 1.031721629e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.3 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.119915666e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.774475196e-08 wvth0 = 1.003084502e-07 pvth0 = -1.252806505e-13
+ k1 = 4.494134777e-01 lk1 = -4.927743860e-08 wk1 = -5.962605746e-07 pk1 = 2.176573958e-12
+ k2 = 2.188907818e-02 lk2 = 2.739723788e-08 wk2 = 2.676290182e-07 pk2 = -9.337719108e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.441809857e-01 ldsub = 6.326443004e-08 wdsub = 1.582317655e-06 pdsub = -6.328107617e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.329197800e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.652705746e-09 wvoff = -9.036340758e-08 pvoff = 4.044496819e-13
+ nfactor = {1.452797052e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.290213634e-07 wnfactor = -3.937492861e-06 pnfactor = 1.516159561e-11
+ eta0 = 7.399584385e-02 leta0 = 2.401221153e-08 weta0 = 6.005735959e-07 peta0 = -2.401852962e-12
+ etab = -6.475108362e-02 letab = -2.099180756e-08 wetab = -5.250297473e-07 petab = 2.099733093e-12
+ u0 = 1.494443245e-02 lu0 = 1.382053321e-11 wu0 = 1.685002563e-08 pu0 = -7.278423250e-14
+ ua = -6.302626519e-10 lua = 2.183945486e-16 wua = 2.554194302e-15 pua = -9.264020289e-21
+ ub = 1.893616172e-18 lub = -3.355714597e-25 wub = -4.943666934e-25 pub = -6.055651387e-31
+ uc = -8.619605630e-11 luc = 3.190362870e-17 wuc = 1.275222280e-16 puc = -2.907828818e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.802866622e+05 lvsat = -2.986430529e-01 wvsat = -6.032978044e-01 pvsat = 1.676987031e-7
+ a0 = 1.121772689e+00 la0 = 1.332043544e-06 wa0 = 5.213475688e-06 pa0 = -1.166125293e-11
+ ags = 1.200413370e-01 lags = 1.095704884e-06 wags = 2.774863816e-06 pags = -3.044017506e-12
+ a1 = 0.0
+ a2 = 1.230120137e+00 la2 = -8.599241350e-07 wa2 = -3.022158278e-06 pa2 = 6.042095269e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.522998383e-02 lketa = -1.808063581e-07 wketa = -6.204490730e-07 pketa = 1.205571483e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.676184906e-01 lpclm = 2.403564029e-06 wpclm = 8.601275643e-06 ppclm = -1.755476015e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 7.234105591e-03 lpdiblc2 = -1.347173793e-08 wpdiblc2 = -4.582507476e-08 ppdiblc2 = 8.807797262e-14
+ pdiblcb = 6.233112532e-04 lpdiblcb = -2.671639850e-09 wpdiblcb = -4.398212555e-09 ppdiblcb = -2.821032770e-15
+ drout = 0.56
+ pscbe1 = 6.848836222e+08 lpscbe1 = 2.301481451e+02 wpscbe1 = 8.088435868e+02 ppscbe1 = -1.617092674e-3
+ pscbe2 = 1.012194425e-08 lpscbe2 = -2.299840379e-15 wpscbe2 = -6.277060888e-15 ppscbe2 = 8.347904324e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.338574203e+00 lbeta0 = 1.656587743e-06 wbeta0 = -7.004714561e-06 pbeta0 = 4.385170507e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.480301510e-11 lagidl = 2.070482588e-16 wagidl = 9.877685154e-16 pagidl = -2.580076494e-21
+ bgidl = 1.332165271e+09 lbgidl = -6.640863996e+02 wbgidl = -2.333896826e+03 pbgidl = 4.666078239e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.276512050e-01 lkt1 = -5.289069037e-08 wkt1 = -3.273614068e-07 pkt1 = 9.837022949e-13
+ kt2 = -3.546941517e-02 lkt2 = -9.243876817e-09 wkt2 = -1.074895902e-08 pkt2 = -2.909414343e-14
+ at = -3.150330841e+05 lat = 1.180583013e+00 wat = 5.263340179e+00 pat = -1.311562777e-5
+ ute = -2.934914571e-01 lute = -2.939708773e-08 wute = -9.580177308e-07 pute = 3.904204437e-12
+ ua1 = 1.929587957e-09 lua1 = 1.065355975e-15 wua1 = 7.530785159e-15 pua1 = -2.386746968e-20
+ ub1 = -5.680795031e-19 lub1 = -8.492323924e-25 wub1 = -5.135803617e-24 pub1 = 1.527367000e-29
+ uc1 = 8.440515145e-11 luc1 = 1.365956172e-16 wuc1 = 1.838595822e-15 puc1 = -6.837123705e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.4 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.099504427e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.062724703e-09 wvth0 = -1.155877452e-07 pvth0 = 3.063530567e-13
+ k1 = 4.209718791e-01 lk1 = 7.584854084e-09 wk1 = 8.719084470e-07 pk1 = -7.586849811e-13
+ k2 = 3.704742328e-02 lk2 = -2.908310938e-09 wk2 = -3.449358634e-07 pk2 = 2.909076172e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.248563615e-01 ldsub = -9.802702512e-08 wdsub = -6.487342653e-06 pdsub = 9.805281799e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.325081924e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.298331457e-10 wvoff = 1.534536107e-07 pvoff = -8.300514914e-14
+ nfactor = {1.307890341e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.068555238e-08 wnfactor = 6.682283711e-06 pnfactor = -6.070151997e-12
+ eta0 = 1.025612777e-01 leta0 = -3.309766049e-08 weta0 = -2.256721398e-06 peta0 = 3.310636915e-12
+ etab = -7.528859417e-02 letab = 7.546846655e-11 wetab = 5.289985705e-07 petab = -7.548832381e-15
+ u0 = 1.487004830e-02 lu0 = 1.625341573e-10 wu0 = -1.142363503e-08 pu0 = -1.625769232e-14
+ ua = -5.150923284e-10 lua = -1.186144832e-17 wua = -2.672965289e-15 pua = 1.186456930e-21
+ ub = 1.701680343e-18 lub = 4.815912575e-26 wub = 1.612214775e-24 pub = -4.817179738e-30
+ uc = -6.957218512e-11 luc = -1.331895119e-18 wuc = -8.455943128e-17 puc = 1.332245567e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.333083536e+05 lvsat = -4.794464738e-03 wvsat = -7.592920936e-01 pvsat = 4.795726258e-7
+ a0 = 1.788772307e+00 la0 = -1.465446683e-09 wa0 = -6.926128788e-07 pa0 = 1.465832272e-13
+ ags = 6.777558291e-01 lags = -1.931417976e-08 wags = 2.859773125e-07 pags = 1.931926170e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.401654004e-02 lketa = -2.378906588e-09 wketa = -1.364620924e-07 pketa = 2.379532526e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.431308069e-01 lpclm = -1.704466486e-08 wpclm = -1.032102182e-06 ppclm = 1.704914966e-12
+ pdiblc1 = 3.865689403e-01 lpdiblc1 = 6.859597592e-09 wpdiblc1 = 3.431962491e-07 ppdiblc1 = -6.861402490e-13
+ pdiblc2 = 5.098128088e-04 lpdiblc2 = -2.809471698e-11 wpdiblc2 = -3.175520202e-09 ppdiblc2 = 2.810210926e-15
+ pdiblcb = -6.979351239e-04 lpdiblcb = -3.011821222e-11 wpdiblcb = -7.316108113e-09 ppdiblcb = 3.012613693e-15
+ drout = 5.818492400e-01 ldrout = -4.368242084e-08 wdrout = -2.185498899e-06 pdrout = 4.369391455e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 9.004194614e-09 lpscbe2 = -6.516264369e-17 wpscbe2 = -5.361761818e-15 ppscbe2 = 6.517978929e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.281925678e+00 lbeta0 = -2.294218441e-07 wbeta0 = 3.450869926e-06 pbeta0 = 2.294822095e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.479667331e-10 lagidl = 7.966481516e-19 wagidl = -2.628864591e-16 pagidl = -7.968577657e-23
+ bgidl = 1.009553072e+09 lbgidl = -1.909912180e+01 wbgidl = -9.555585256e+02 pbgidl = 1.910414716e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.571418188e-01 lkt1 = 6.068861640e-09 wkt1 = 4.683050720e-07 pkt1 = -6.070458479e-13
+ kt2 = -4.035669769e-02 lkt2 = 5.270960712e-10 wkt2 = 1.070050789e-09 pkt2 = -5.272347607e-14
+ at = 2.796664617e+05 lat = -8.378974042e-03 wat = -1.716097587e+00 pat = 8.381178718e-7
+ ute = -4.021138694e-01 lute = 1.877678994e-07 wute = 1.038911980e-05 pute = -1.878173049e-11
+ ua1 = 2.275221051e-09 lua1 = 3.743438287e-16 wua1 = 1.432166227e-14 pua1 = -3.744423260e-20
+ ub1 = -8.870950591e-19 lub1 = -2.114357569e-25 wub1 = -8.074618125e-24 pub1 = 2.114913898e-29
+ uc1 = 1.581694808e-10 luc1 = -1.087882474e-17 wuc1 = -2.125507197e-15 puc1 = 1.088168717e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.5 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.106160919e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.588875093e-09 wvth0 = 5.270001767e-08 pvth0 = 1.381889853e-13
+ k1 = 3.612078053e-01 lk1 = 6.730500130e-08 wk1 = 3.417309195e-07 pk1 = -2.288971340e-13
+ k2 = 6.167805224e-02 lk2 = -2.752083639e-08 wk2 = -1.728979393e-07 pk2 = 1.189961411e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.517077494e-01 ldsub = -2.247851772e-07 wdsub = 1.744578820e-06 pdsub = 1.579410788e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.472361426e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.554695826e-08 wvoff = 1.472363370e-07 pvoff = -7.679244517e-14
+ nfactor = {9.127602572e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.555252152e-07 wnfactor = -1.982904471e-06 pnfactor = 2.588667272e-12
+ eta0 = 1.393095928e-01 leta0 = -6.981896560e-08 weta0 = 2.007882397e-06 peta0 = -9.508323971e-13
+ etab = -1.498540325e-01 letab = 7.458610121e-08 wetab = 1.045894875e-06 petab = -5.240652180e-13
+ u0 = 1.761672575e-02 lu0 = -2.582124484e-09 wu0 = -2.770868176e-08 pu0 = 1.538489589e-17
+ ua = -2.471997206e-10 lua = -2.795571550e-16 wua = -1.985304443e-15 pua = 4.993015152e-22
+ ub = 1.845505706e-18 lub = -9.556052554e-26 wub = -2.237107196e-24 pub = -9.706870189e-31
+ uc = -6.465566351e-11 luc = -6.244803083e-18 wuc = -3.394659725e-16 puc = 3.879437416e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.995301843e+05 lvsat = -7.096762239e-02 wvsat = -5.183317586e-01 pvsat = 2.387893966e-7
+ a0 = 1.828111619e+00 la0 = -4.077584408e-08 wa0 = 3.557327537e-06 pa0 = -4.100233482e-12
+ ags = 4.775075328e-01 lags = 1.807869341e-07 wags = 3.765105471e-06 pags = -1.544644829e-12
+ a1 = 0.0
+ a2 = 8.150873818e-01 la2 = -1.507629254e-08 wa2 = -1.509135156e-06 pa2 = 1.508025942e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.307606676e-02 lketa = -3.318688619e-09 wketa = -1.549988315e-11 pketa = 1.016069483e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.641678557e-01 lpclm = -3.806625144e-08 wpclm = -7.662274314e-07 ppclm = 1.439235633e-12
+ pdiblc1 = 3.716491251e-01 lpdiblc1 = 2.176844674e-08 wpdiblc1 = 1.835570341e-06 ppdiblc1 = -2.177417446e-12
+ pdiblc2 = 7.593741736e-04 lpdiblc2 = -2.774726542e-10 wpdiblc2 = -4.746354507e-09 ppdiblc2 = 4.379890668e-15
+ pdiblcb = -1.687414322e-03 lpdiblcb = 9.586337183e-10 wpdiblcb = 1.684357973e-07 ppdiblcb = -1.726101141e-13
+ drout = 5.459672928e-01 ldrout = -7.826846833e-09 wdrout = 1.403639951e-06 pdrout = 7.828906233e-13
+ pscbe1 = 7.969043332e+08 lpscbe1 = 3.093391532e+00 wpscbe1 = 3.096481379e+02 ppscbe1 = -3.094205465e-4
+ pscbe2 = 9.239998590e-09 lpscbe2 = -3.007933040e-16 wpscbe2 = -1.172896844e-15 ppscbe2 = 2.332192771e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.950169287e+00 lbeta0 = 2.100620706e-06 wbeta0 = 3.937602814e-05 pbeta0 = -1.295053227e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.917878126e-10 lagidl = -4.299222289e-17 wagidl = -6.449298092e-16 pagidl = 3.020767716e-22
+ bgidl = 9.936517962e+08 lbgidl = -3.209533790e+00 wbgidl = 6.349874132e+02 pbgidl = 3.210378282e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.759413225e-01 lkt1 = 2.485454764e-08 wkt1 = 1.723807220e-07 pkt1 = -3.113390023e-13
+ kt2 = -3.513807962e-02 lkt2 = -4.687686320e-09 wkt2 = -1.865332619e-07 pkt2 = 1.347419482e-13
+ at = 4.475575579e+05 lat = -1.761466703e-01 wat = -1.369342664e+00 pat = 4.916178143e-7
+ ute = -2.574618304e-01 lute = 4.322217970e-08 wute = -1.722769808e-05 pute = 8.814789031e-12
+ ua1 = 3.518452698e-09 lua1 = -8.679740430e-16 wua1 = -5.178462214e-14 pua1 = 2.861346368e-20
+ ub1 = -1.669408731e-18 lub1 = 5.703029144e-25 wub1 = 3.708533246e-23 pub1 = -2.397761903e-29
+ uc1 = 3.572772385e-10 luc1 = -2.098402383e-16 wuc1 = -1.143282140e-15 puc1 = 1.066655951e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.6 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.099385702e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.062464225e-10 wvth0 = 3.708057417e-07 pvth0 = -2.063006900e-14
+ k1 = 5.161882560e-01 lk1 = -1.007131342e-08 wk1 = -2.134496079e-06 pk1 = 1.007396339e-12
+ k2 = -3.228630546e-04 lk2 = 3.434050585e-09 wk2 = 7.534469003e-07 pk2 = -3.434954153e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.776351188e-01 ldsub = 1.190269470e-08 wdsub = 7.292721473e-06 pdsub = -1.190582654e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.184110015e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.155574195e-09 wvoff = 2.249413230e-07 pvoff = -1.155878250e-13
+ nfactor = {1.806697789e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.213493560e-09 wnfactor = 5.047948991e-06 pnfactor = -9.215917815e-13
+ eta0 = 3.530907186e-02 leta0 = -1.789514552e-08 weta0 = -3.481823083e-06 peta0 = 1.789985409e-12
+ etab = -4.339755216e-04 letab = -1.410354099e-11 wetab = -6.604185076e-09 petab = 1.410725191e-15
+ u0 = 1.218175985e-02 lu0 = 1.313637656e-10 wu0 = -1.359512679e-09 pu0 = -1.313983301e-14
+ ua = -8.779859040e-10 lua = 3.537230888e-17 wua = 6.101509411e-15 pua = -3.538161604e-21
+ ub = 1.704935269e-18 lub = -2.537862623e-26 wub = -9.265874293e-24 pub = 2.538530386e-30
+ uc = -7.604056516e-11 luc = -5.607201649e-19 wuc = 3.252250662e-16 puc = 5.608677016e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.971604343e+04 lvsat = -1.163315347e-03 wvsat = -2.731167869e-01 pvsat = 1.163621438e-7
+ a0 = 1.723694094e+00 la0 = 1.135617120e-08 wa0 = -2.380035503e-06 pa0 = -1.135915924e-12
+ ags = 9.428943723e-01 lags = -5.156442633e-08 wags = -9.659517174e-06 pags = 5.157799396e-12
+ a1 = 0.0
+ a2 = 7.698252365e-01 la2 = 7.521512433e-09 wa2 = 3.018270312e-06 pa2 = -7.523491493e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.399726728e-02 lketa = 2.133884556e-09 wketa = 6.310152167e-07 pketa = -2.134446024e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.753450874e-01 lpclm = 6.279847967e-09 wpclm = 3.374630961e-06 ppclm = -6.281500321e-13
+ pdiblc1 = 4.392819450e-01 lpdiblc1 = -1.199825307e-08 wpdiblc1 = -4.929491202e-06 ppdiblc1 = 1.200141005e-12
+ pdiblc2 = 7.832012369e-04 lpdiblc2 = -2.893686730e-10 wpdiblc2 = -5.394786172e-08 ppdiblc2 = 2.894448117e-14
+ pdiblcb = 2.326756472e-04 wpdiblcb = -1.772926517e-7
+ drout = 5.008305208e-01 ldrout = 1.470836363e-08 wdrout = 5.918504788e-06 pdrout = -1.471223370e-12
+ pscbe1 = 8.061913337e+08 lpscbe1 = -1.543282793e+00 wpscbe1 = -6.192962758e+02 ppscbe1 = 1.543688862e-4
+ pscbe2 = 8.024688260e-09 lpscbe2 = 3.059686081e-16 wpscbe2 = 6.479828924e-14 ppscbe2 = -3.060491145e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.281234578e-09 lalpha0 = -5.897490816e-16 walpha0 = -1.181545385e-13 palpha0 = 5.899042564e-20
+ alpha1 = 9.246703802e-11 lalpha1 = 3.760944264e-18 walpha1 = 7.534944054e-16 palpha1 = -3.761933843e-22
+ beta0 = 7.728521072e+00 lbeta0 = -2.850430978e-07 wbeta0 = -4.367073480e-05 pbeta0 = 2.851180983e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.056767836e-10 wagidl = -3.988685277e-17
+ bgidl = 9.927359681e+08 lbgidl = -2.752292861e+00 wbgidl = 7.265943230e+02 pbgidl = 2.753017044e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.266494521e-01 lkt1 = 2.448419847e-10 wkt1 = -4.021605767e-07 pkt1 = -2.449064075e-14
+ kt2 = -4.495712659e-02 lkt2 = 2.146201649e-10 wkt2 = 1.263458940e-07 pkt2 = -2.146766357e-14
+ at = 9.514384745e+04 lat = -1.988391675e-04 wat = -4.244964088e-01 pat = 1.988914861e-8
+ ute = -1.663704336e-01 lute = -2.256566558e-09 wute = -2.426302467e-08 pute = 2.257160306e-13
+ ua1 = 1.677240366e-09 lua1 = 5.127883150e-17 wua1 = 1.580011959e-14 pua1 = -5.129232399e-21
+ ub1 = -4.260849844e-19 lub1 = -5.044511591e-26 wub1 = -2.104703800e-23 pub1 = 5.045838903e-30
+ uc1 = -5.389193781e-11 luc1 = -4.557859431e-18 wuc1 = -1.842790967e-15 puc1 = 4.559058695e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.7 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.110990219e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.098846321e-09 wvth0 = 1.531562767e-06 pvth0 = -3.099661689e-13
+ k1 = 5.216229468e-01 lk1 = -1.142599163e-08 wk1 = -2.678108160e-06 pk1 = 1.142899804e-12
+ k2 = -3.258953263e-03 lk2 = 4.165915111e-09 wk2 = 1.047133176e-06 pk2 = -4.167011247e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.024539681e-01 ldsub = 5.716224228e-09 wdsub = 4.810183509e-06 pdsub = -5.717728281e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.196347135e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.460602765e-09 wvoff = 3.473447204e-07 pvoff = -1.460987078e-13
+ nfactor = {1.834543320e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.272577329e-09 wnfactor = 2.262663241e-06 pnfactor = -2.273175289e-13
+ eta0 = -3.648257768e-02 weta0 = 3.699230853e-6
+ etab = -4.905560381e-04 letab = 1.446853325e-18 wetab = -9.446446833e-10 petab = -1.447234012e-22
+ u0 = 1.236528989e-02 lu0 = 8.561615126e-11 wu0 = -1.971734530e-08 pu0 = -8.563867858e-15
+ ua = -8.091883400e-10 lua = 1.822348407e-17 wua = -7.800571972e-16 pua = -1.822827903e-21
+ ub = 1.636971215e-18 lub = -8.437566263e-27 wub = -2.467680602e-24 pub = 8.439786355e-31
+ uc = -8.041065455e-11 luc = 5.285901684e-19 wuc = 7.623489917e-16 puc = -5.287292511e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.562071131e+04 lvsat = -1.424923844e-04 wvsat = 1.365241820e-01 pvsat = 1.425298770e-8
+ a0 = 1.735006299e+00 la0 = 8.536434573e-09 wa0 = -3.511553590e-06 pa0 = -8.538680679e-13
+ ags = 5.316721438e-01 lags = 5.093888246e-08 wags = 3.147352576e-05 pags = -5.095228550e-12
+ a1 = 0.0
+ a2 = 7.854091278e-01 la2 = 3.636993767e-09 wa2 = 1.459471138e-06 pa2 = -3.637950733e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.557528761e-02 lketa = 3.457979429e-11 wketa = -2.114043492e-07 pketa = -3.458889292e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.968691212e-01 lpclm = 9.146596731e-10 wpclm = 1.221661237e-06 ppclm = -9.149003384e-14
+ pdiblc1 = 3.974874942e-01 lpdiblc1 = -1.580359296e-09 wpdiblc1 = -7.489464268e-07 ppdiblc1 = 1.580775120e-13
+ pdiblc2 = -2.488458694e-04 lpdiblc2 = -3.211545102e-11 wpdiblc2 = 4.928400414e-08 ppdiblc2 = 3.212390124e-15
+ pdiblcb = -2.886522699e-02 lpdiblcb = 7.253088702e-09 wpdiblcb = 2.733263236e-06 ppdiblcb = -7.254997135e-13
+ drout = 5.642746893e-01 ldrout = -1.106047019e-09 wdrout = -4.275814013e-07 pdrout = 1.106338042e-13
+ pscbe1 = 7.999802145e+08 lpscbe1 = 4.931840675e-03 wpscbe1 = 1.979073813e+00 ppscbe1 = -4.933138341e-7
+ pscbe2 = 1.085463318e-08 lpscbe2 = -3.994376134e-16 wpscbe2 = -2.182706646e-13 ppscbe2 = 3.995427134e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.330249408e-09 lalpha0 = 6.120247407e-17 walpha0 = 1.430625735e-13 palpha0 = -6.121857766e-21
+ alpha1 = 1.075551742e-10 walpha1 = -7.557162111e-16
+ beta0 = 6.495175930e+00 lbeta0 = 2.238667910e-08 wbeta0 = 7.969623120e-05 pbeta0 = -2.239256948e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.056767836e-10 wagidl = -3.988685277e-17
+ bgidl = 1.011677155e+09 lbgidl = -7.473667760e+00 wbgidl = -1.168022726e+03 pbgidl = 7.475634231e-4
+ cgidl = 2.514436011e+02 lcgidl = 1.210341077e-05 wcgidl = 4.856917504e-03 pcgidl = -1.210659542e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.296922307e-01 lkt1 = 1.003300177e-09 wkt1 = -9.780266133e-08 pkt1 = -1.003564165e-13
+ kt2 = -4.694308991e-02 lkt2 = 7.096513130e-10 wkt2 = 3.249944811e-07 pkt2 = -7.098380364e-14
+ at = 9.197425222e+04 lat = 5.912299861e-04 wat = -1.074534880e-01 pat = -5.913855505e-8
+ ute = -1.980491722e-01 lute = 5.639834231e-09 wute = 3.144444371e-06 pute = -5.641318185e-13
+ ua1 = 1.723253439e-09 lua1 = 3.980938291e-17 wua1 = 1.119760161e-14 pua1 = -3.981985755e-21
+ ub1 = -4.710933944e-19 lub1 = -3.922609460e-26 wub1 = -1.654501274e-23 pub1 = 3.923641577e-30
+ uc1 = -5.964273257e-11 luc1 = -3.124387574e-18 wuc1 = -1.267560175e-15 puc1 = 3.125209663e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.8 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-1.103484708e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.919646093e-09 wvth0 = 7.808142354e-07 pvth0 = -1.920151190e-13
+ k1 = 4.989864323e-01 lk1 = -8.066782026e-09 wk1 = -4.138610987e-07 pk1 = 8.068904557e-13
+ k2 = -8.790807193e-03 lk2 = 5.646685125e-09 wk2 = 1.600464123e-06 pk2 = -5.648170881e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.272539581e-01 ldsub = 2.101743331e-08 wdsub = 1.233216318e-05 pdsub = -2.102296342e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.262644455e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.900298519e-09 wvoff = 1.010492361e-06 pvoff = -2.901061646e-13
+ nfactor = {2.259544656e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.092479758e-08 wnfactor = -4.024865300e-05 pnfactor = 8.094609052e-12
+ eta0 = -1.495370710e-01 leta0 = 2.218864014e-08 weta0 = 1.500765488e-05 peta0 = -2.219447841e-12
+ etab = -1.524171035e-02 letab = 2.895135303e-09 wetab = 1.474558919e-06 petab = -2.895897071e-13
+ u0 = 1.345813674e-02 lu0 = -1.207523136e-10 wu0 = -1.290307857e-07 pu0 = 1.207840860e-14
+ ua = -5.043885668e-10 lua = -3.986987992e-17 wua = -3.126805441e-14 pua = 3.988037048e-21
+ ub = 1.399444518e-18 lub = 3.738046242e-26 wub = 2.129123891e-23 pub = -3.739029797e-30
+ uc = -7.916584896e-11 luc = 3.344054886e-19 wuc = 6.378356788e-16 puc = -3.344934774e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.735587026e+04 lvsat = 1.466093852e-03 wvsat = 9.632257510e-01 pvsat = -1.466479611e-7
+ a0 = 1.777625859e+00 la0 = 9.812309750e-10 wa0 = -7.774631013e-06 pa0 = -9.814891565e-14
+ ags = 8.158262311e-01 wags = 3.050640362e-6
+ a1 = 0.0
+ a2 = 8.305062086e-01 la2 = -4.869082588e-09 wa2 = -3.051423535e-06 pa2 = 4.870363741e-13
+ b0 = 8.823693846e-25 lb0 = -1.731782273e-31 wb0 = -8.826015537e-29 pb0 = 1.732237939e-35
+ b1 = 0.0
+ keta = -2.752911257e-02 lketa = -5.466623489e-09 wketa = -3.016759804e-06 pketa = 5.468061867e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.704227881e-01 lpclm = 6.191887955e-09 wpclm = 3.866990407e-06 ppclm = -6.193517164e-13
+ pdiblc1 = 2.927906757e-01 lpdiblc1 = 1.881809366e-08 wpdiblc1 = 9.723490201e-06 ppdiblc1 = -1.882304508e-12
+ pdiblc2 = -2.638915872e-03 lpdiblc2 = 4.339260760e-10 wpdiblc2 = 2.883538919e-07 ppdiblc2 = -4.340402506e-14
+ pdiblcb = 1.437533867e-02 lpdiblcb = -5.456983758e-10 wpdiblcb = -1.591931075e-06 ppdiblcb = 5.458419599e-14
+ drout = 7.318381714e-01 ldrout = -3.409778213e-08 wdrout = -1.718833855e-05 pdrout = 3.410675394e-12
+ pscbe1 = 8.000505443e+08 lpscbe1 = -8.403742002e-03 wpscbe1 = -5.055756289e+00 ppscbe1 = 8.405953195e-7
+ pscbe2 = 8.723860191e-09 lpscbe2 = -1.912078944e-17 wpscbe2 = -5.137300497e-15 ppscbe2 = 1.912582051e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -4.706165106e-09 lalpha0 = 7.295805016e-16 walpha0 = 4.807429704e-13 palpha0 = -7.297724689e-20
+ alpha1 = 1.075551742e-10 walpha1 = -7.557162111e-16
+ beta0 = 5.641366997e+00 lbeta0 = 1.920824556e-07 wbeta0 = 1.650995899e-04 pbeta0 = -1.921329963e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.056767836e-10 wagidl = -3.988685277e-17
+ bgidl = 9.226506253e+08 lbgidl = 9.290383626e+00 wbgidl = 7.736972688e+03 pbgidl = -9.292828112e-4
+ cgidl = 4.240425281e+02 lcgidl = -2.062393093e-05 wcgidl = -1.240751661e-02 pcgidl = 2.062935750e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.286386032e-01 lkt1 = 8.916546130e-10 wkt1 = -2.031931333e-07 pkt1 = -8.918892251e-14
+ kt2 = -3.774706395e-02 lkt2 = -1.027909299e-09 wkt2 = -5.948500803e-07 pkt2 = 1.028179763e-13
+ at = 9.182333092e+04 lat = 6.769178845e-04 wat = -9.235738681e-02 pat = -6.770959952e-8
+ ute = -2.139288169e-01 lute = 9.291287608e-09 wute = 4.732826661e-06 pute = -9.293732331e-13
+ ua1 = 1.960095917e-09 lua1 = -2.899315645e-18 wua1 = -1.249287799e-14 pua1 = 2.900078513e-22
+ ub1 = -7.368343748e-19 lub1 = 9.209682720e-27 wub1 = 1.003607748e-23 pub1 = -9.212105972e-31
+ uc1 = -8.847851451e-11 luc1 = 2.238776264e-18 wuc1 = 1.616776745e-15 puc1 = -2.239365331e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.9 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.104325265e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.462794766e-07 wvth0 = -3.838358253e-08 pvth0 = 3.838330041e-12
+ k1 = 4.350683671e-01 lk1 = 1.503441838e-07 wk1 = 1.056372907e-08 pk1 = -1.056365143e-12
+ k2 = 3.092240711e-02 lk2 = -1.841405577e-07 wk2 = -1.293838520e-08 pk2 = 1.293829010e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.337777855e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.378895320e-07 wvoff = 9.688619944e-09 pvoff = -9.688548732e-13
+ nfactor = {1.389953464e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.114106249e-07 wnfactor = 2.890720657e-08 pnfactor = -2.890699410e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.416129041e-02 lu0 = 7.731019075e-08 wu0 = 5.432095136e-09 pu0 = -5.432055210e-13
+ ua = -5.198134195e-10 lua = -5.346315750e-15 wua = -3.756515861e-16 pua = 3.756488251e-20
+ ub = 1.608654607e-18 lub = 1.945956926e-23 wub = 1.367300100e-24 pub = -1.367290050e-28
+ uc = -7.885570791e-11 luc = 1.185003204e-16 wuc = 8.326263434e-18 puc = -8.326202236e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.750656967e+05 lvsat = 2.493412005e+00 wvsat = 1.751961946e-01 pvsat = -1.751949069e-5
+ a0 = 1.585351506e+00 la0 = -1.075357159e-05 wa0 = -7.555850445e-07 pa0 = 7.555794910e-11
+ ags = 5.006254759e-01 lags = -8.647504032e-06 wags = -6.076050794e-07 pags = 6.076006135e-11
+ a1 = 0.0
+ a2 = 8.743431006e-01 la2 = 1.256459759e-05 wa2 = 8.828343171e-07 pa2 = -8.828278283e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.636629039e-02 lketa = 2.319703789e-06 wketa = 1.629908237e-07 pketa = -1.629896257e-11
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.382975169e-01 lpclm = -6.280739325e-06 wpclm = -4.413075845e-07 ppclm = 4.413043409e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.453037867e-03 lpdiblc2 = 2.174545550e-07 wpdiblc2 = 1.527914780e-08 ppdiblc2 = -1.527903549e-12
+ pdiblcb = -1.961401813e-03 lpdiblcb = 1.865644062e-07 wpdiblcb = 1.310869361e-08 ppdiblcb = -1.310859726e-12
+ drout = 0.56
+ pscbe1 = 7.290520221e+08 lpscbe1 = 1.742297986e+03 wpscbe1 = 1.224201923e+02 ppscbe1 = -1.224192925e-2
+ pscbe2 = 9.567772474e-09 lpscbe2 = -6.277951227e-15 wpscbe2 = -4.411116826e-16 ppscbe2 = 4.411084404e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.353153947e-10 lalpha0 = -2.353136651e-14 walpha0 = -1.653399381e-15 palpha0 = 1.653387229e-19
+ alpha1 = 3.734635130e-11 lalpha1 = 6.265318820e-15 walpha1 = 4.402240837e-16 palpha1 = -4.402208481e-20
+ beta0 = 3.801232528e+00 lbeta0 = 9.911492874e-05 wbeta0 = 6.964175319e-06 pbeta0 = -6.964124132e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.340389132e+09 lbgidl = -1.859431650e+04 wbgidl = -1.306504294e+03 pbgidl = 1.306494692e-1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.354073409e-01 lkt1 = -6.282612926e-07 wkt1 = -4.414392305e-08 pkt1 = 4.414359860e-12
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.321172741e-01 lute = 3.145704292e-06 wute = 2.210286227e-07 pute = -2.210269982e-11
+ ua1 = 2.2116e-9
+ ub1 = -8.733609226e-19 lub1 = 7.977033632e-24 wub1 = 5.604953910e-25 pub1 = -5.604912714e-29
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.10 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.131640243e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.535399727e-7
+ k1 = 4.425858526e-01 wk1 = -4.225646922e-8
+ k2 = 2.171504086e-02 wk2 = 5.175544281e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.268830555e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff = -3.875590405e-8
+ nfactor = {1.410524751e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.156330758e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.802694201e-02 wu0 = -2.172917909e-8
+ ua = -7.871390313e-10 wua = 1.502661567e-15
+ ub = 2.581668828e-18 wub = -5.469401399e-24
+ uc = -7.293047414e-11 wuc = -3.330627774e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.997408787e+05 wvsat = -7.008105333e-1
+ a0 = 1.047653166e+00 wa0 = 3.022451253e-6
+ ags = 6.823438395e-02 wags = 2.430509639e-6
+ a1 = 0.0
+ a2 = 1.502596068e+00 wa2 = -3.531467050e-6
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.962316167e-02 wketa = -6.519872552e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.757509907e-01 wpclm = 1.765295213e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.232616521e-02 wpdiblc2 = -6.111883730e-8
+ pdiblcb = 7.367161319e-03 wpdiblcb = -5.243670147e-8
+ drout = 0.56
+ pscbe1 = 8.161701230e+08 wpscbe1 = -4.896987655e+2
+ pscbe2 = 9.253863376e-09 wpscbe2 = 1.764511576e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.412961713e-10 walpha0 = 6.613840584e-15
+ alpha1 = 3.506238052e-10 walpha1 = -1.760961050e-15
+ beta0 = 8.757161095e+00 wbeta0 = -2.785772505e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 4.106391384e+08 wbgidl = 5.226209240e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.668215600e-01 wkt1 = 1.765821816e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -1.748262791e-01 wute = -8.841469833e-7
+ ua1 = 2.2116e-9
+ ub1 = -4.744945827e-19 wub1 = -2.242063960e-24
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.11 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.146089557e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.155838927e-07 wvth0 = 1.909402685e-07 pvth0 = -2.991748771e-13
+ k1 = 6.149778499e-01 lk1 = -1.379009271e-06 wk1 = -1.205182156e-06 pk1 = 9.302550745e-12
+ k2 = -5.102097423e-02 lk2 = 5.818346597e-07 wk2 = 5.310824463e-07 pk2 = -3.834263723e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.454280064e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.483459769e-07 wvoff = 8.153731693e-08 pvoff = -9.622573524e-13
+ nfactor = {1.027096500e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.067144186e-06 wnfactor = 2.714542149e-06 pnfactor = -2.263932162e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.547945506e-02 lu0 = 2.037802316e-08 wu0 = -2.575381360e-09 pu0 = -1.532163038e-13
+ ua = -1.246522019e-09 lua = 3.674726256e-15 wua = 4.509408419e-15 pua = -2.405176485e-20
+ ub = 2.722066113e-18 lub = -1.123075088e-24 wub = -5.855564044e-24 pub = 3.089017325e-30
+ uc = -1.289533508e-10 luc = 4.481418365e-16 wuc = 3.093744797e-16 puc = -2.741194189e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.976226949e+05 lvsat = -7.829825860e-01 wvsat = -8.667221047e-01 pvsat = 1.327170627e-6
+ a0 = 2.075952360e-01 la0 = 6.719846001e-06 wa0 = 6.789122187e-06 pa0 = -3.013059896e-11
+ ags = -5.949870005e-01 lags = 5.305283608e-06 wags = 5.218587462e-06 pags = -2.230257335e-11
+ a1 = 0.0
+ a2 = 2.205063035e+00 la2 = -5.619219418e-06 wa2 = -7.062285193e-06 pa2 = 2.824394999e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.241315780e-01 lketa = -1.155961117e-06 wketa = -1.370810259e-06 pketa = 5.750055695e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -9.841659078e-01 lpclm = 6.466725152e-06 wpclm = 3.530266052e-06 ppclm = -1.411846946e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 2.351108305e-02 lpdiblc2 = -8.947112183e-08 wpdiblc2 = -1.175820215e-07 ppdiblc2 = 4.516639729e-13
+ pdiblcb = 9.775365094e-03 lpdiblcb = -1.926386016e-08 wpdiblcb = -6.461326466e-08 ppdiblcb = 9.740355569e-14
+ drout = 0.56
+ pscbe1 = 6.413643235e+08 lpscbe1 = 1.398317913e+03 wpscbe1 = 3.625279895e+02 ppscbe1 = -6.817187654e-3
+ pscbe2 = 9.814620529e-09 lpscbe2 = -4.485645066e-15 wpscbe2 = 1.719138294e-15 ppscbe2 = 3.629529050e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.782419379e-09 lalpha0 = 7.528293939e-15 walpha0 = 1.322646587e-14 palpha0 = -5.289614204e-20
+ alpha1 = 6.012015583e-10 lalpha1 = -2.004437850e-15 walpha1 = -3.521598524e-15 palpha1 = 1.408380572e-20
+ beta0 = 1.383573023e+01 lbeta0 = -4.062482035e-05 wbeta0 = -6.722270159e-05 pbeta0 = 3.148908791e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 9.349118961e-09 lagidl = -7.398615359e-14 wagidl = -6.530569988e-14 pagidl = 5.223975993e-19
+ bgidl = 2.401991617e+09 lbgidl = -1.592935619e+04 wbgidl = -7.680678031e+03 pbgidl = 1.032456116e-1
+ cgidl = 300.0
+ egidl = 6.271194736e-01 legidl = -4.216568356e-06 wegidl = -3.703705883e-06 pegidl = 2.962692484e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.389169645e-01 lkt1 = -2.232162542e-07 wkt1 = 5.617526259e-08 pkt1 = 9.631668531e-13
+ kt2 = -4.614231739e-02 lkt2 = 6.544452582e-08 wkt2 = 7.423916341e-08 pkt2 = -5.938587415e-13
+ at = -4.620701916e+05 lat = 3.696221912e+00 wat = 1.402511092e+00 pat = -1.121905789e-5
+ ute = -2.297145685e+00 lute = 1.697699534e-05 wute = 1.401100103e-05 pute = -1.191502362e-10
+ ua1 = -4.920624649e-09 lua1 = 5.705255500e-14 wua1 = 4.866046131e-14 pua1 = -3.892479250e-19
+ ub1 = 4.319015307e-18 lub1 = -3.834455589e-23 wub1 = -3.469879062e-23 pub1 = 2.596299576e-28
+ uc1 = -8.888517754e-11 luc1 = 1.669728000e-15 wuc1 = 1.346721376e-15 puc1 = -1.077278117e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.12 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.117839253e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.603443242e-09 wvth0 = 8.571892767e-08 pvth0 = 1.216331486e-13
+ k1 = 1.425366097e-01 lk1 = 5.104084460e-07 wk1 = 1.559952046e-06 pk1 = -1.755953689e-12
+ k2 = 1.501357501e-01 lk2 = -2.226443875e-07 wk2 = -6.334721118e-07 pk2 = 8.230985621e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.295584163e+00 ldsub = -2.941795997e-06 wdsub = -3.697275504e-06 pdsub = 1.478638452e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.417604178e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.336783184e-07 wvoff = -2.824632783e-08 pvoff = -5.232034643e-13
+ nfactor = {1.687630973e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.499846922e-06 wnfactor = 5.084530321e-06 pnfactor = -3.211753237e-11
+ eta0 = 3.591932608e-01 leta0 = -1.116567836e-06 weta0 = -1.403312437e-06 peta0 = 5.612218313e-12
+ etab = -3.140746116e-01 letab = 9.761190516e-07 wetab = 1.226795149e-06 petab = -4.906278902e-12
+ u0 = 2.285056832e-02 lu0 = -9.101012085e-09 wu0 = -3.870095171e-08 pu0 = -8.740574691e-15
+ ua = -4.061905855e-10 lua = 3.140181655e-16 wua = 9.797940533e-16 pua = -9.935901656e-21
+ ub = 2.949120190e-18 lub = -2.031124510e-24 wub = -7.910667240e-24 pub = 1.130791961e-29
+ uc = 7.121539226e-11 luc = -3.523860117e-16 wuc = -9.784997220e-16 puc = 2.409356030e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.929805420e+05 lvsat = -3.644908864e-01 wvsat = -6.924889641e-01 pvsat = 6.303661257e-7
+ a0 = 1.915628181e+00 la0 = -1.110303737e-07 wa0 = -3.644006768e-07 pa0 = -1.521765349e-12
+ ags = 6.963522212e-01 lags = 1.408758555e-07 wags = -1.274476265e-06 pags = 3.664909157e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.728837900e-02 lketa = 8.948981748e-08 wketa = 2.404031700e-07 pketa = -6.936137789e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.731781465e-01 lpclm = 1.438273083e-06 wpclm = 2.693576142e-06 ppclm = -1.077232479e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.961675541e-03 lpdiblc2 = -3.289330615e-09 wpdiblc2 = -8.779336231e-09 ppdiblc2 = 1.653320194e-14
+ pdiblcb = 1.144856022e-02 lpdiblcb = -2.595541089e-08 wpdiblcb = -8.045978931e-08 ppdiblcb = 1.607780071e-13
+ drout = 0.56
+ pscbe1 = 1.180613741e+09 lpscbe1 = -7.582834076e+02 wpscbe1 = -2.674310895e+03 ppscbe1 = 5.327935806e-3
+ pscbe2 = 9.695501107e-09 lpscbe2 = -4.009254933e-15 wpscbe2 = -3.280738287e-15 ppscbe2 = 2.035878432e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.784652466e-03 lalpha0 = -1.113656275e-08 walpha0 = -1.956583634e-08 palpha0 = 7.824896446e-14
+ alpha1 = -1.512232415e-10 lalpha1 = 1.004708317e-15 walpha1 = 1.765172877e-15 palpha1 = -7.059394104e-21
+ beta0 = 6.785632980e+01 lbeta0 = -2.566675135e-04 wbeta0 = -4.533002829e-04 pbeta0 = 1.858917437e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.841677362e-08 lagidl = 3.705700879e-14 wagidl = 1.307045659e-13 pagidl = -2.614993964e-19
+ bgidl = -3.321663720e+09 lbgidl = 6.961058278e+03 wbgidl = 3.036535766e+04 pbgidl = -4.891056731e-2
+ cgidl = 300.0
+ egidl = -9.542389472e-01 legidl = 2.107703029e-06 wegidl = 7.407411766e-06 pegidl = -1.480937908e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.882970012e-01 lkt1 = 3.741940984e-07 wkt1 = 8.013860787e-07 pkt1 = -2.017128681e-12
+ kt2 = -2.946525915e-02 lkt2 = -1.251449469e-09 wkt2 = -5.293603250e-08 pkt2 = -8.525143161e-14
+ at = 7.381904975e+05 lat = -1.103938654e+00 wat = -2.136937312e+00 pat = 2.936134230e-6
+ ute = 4.310534268e+00 lute = -9.448867823e-06 wute = -3.330733893e-05 pute = 7.008834469e-11
+ ua1 = 1.785963804e-08 lua1 = -3.405175225e-14 wua1 = -1.043987169e-13 pua1 = 2.228762892e-19
+ ub1 = -1.146452347e-17 lub1 = 2.477799831e-23 wub1 = 7.142601138e-23 pub1 = -1.647912486e-28
+ uc1 = 1.048320467e-09 luc1 = -2.878258730e-15 wuc1 = -4.934173924e-15 puc1 = 1.434618358e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.13 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.153718427e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.433541902e-08 wvth0 = 2.653367362e-07 pvth0 = -2.374704493e-13
+ k1 = 3.428299086e-01 lk1 = 1.099690637e-07 wk1 = 1.420958312e-06 pk1 = -1.478068381e-12
+ k2 = 4.790378036e-02 lk2 = -1.825558849e-08 wk2 = -4.212160155e-07 pk2 = 3.987423777e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.719093182e+00 ldsub = 3.085342905e-06 wdsub = 9.981978152e-06 pdsub = -1.256206854e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.317410751e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.627950286e-08 wvoff = -5.545675949e-07 pvoff = 5.290522237e-13
+ nfactor = {5.927061865e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.012518263e-06 wnfactor = -2.577345660e-05 pnfactor = 2.957576085e-11
+ eta0 = -6.175161750e-01 leta0 = 8.361331540e-07 weta0 = 2.802767448e-06 peta0 = -2.796849988e-12
+ etab = -4.108820591e-01 letab = 1.169662793e-06 wetab = 2.886982960e-06 petab = -8.225434287e-12
+ u0 = 2.380166608e-02 lu0 = -1.100250854e-08 wu0 = -7.417996818e-08 pu0 = 6.219138117e-14
+ ua = 4.188241201e-10 lua = -1.335404860e-15 wua = -9.234953638e-15 pua = 1.048608589e-20
+ ub = 2.031643100e-18 lub = -1.968446761e-25 wub = -7.062065040e-25 pub = -3.095706585e-30
+ uc = -1.278323047e-10 luc = 4.556308219e-17 wuc = 3.247943462e-16 puc = -1.962741851e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.228770102e+04 lvsat = 3.674728633e-02 wvsat = -4.710681900e-01 pvsat = 1.876873218e-7
+ a0 = 5.941576999e-01 la0 = 2.530939307e-06 wa0 = 7.701122070e-06 pa0 = -1.764688268e-11
+ ags = -4.032361232e-01 lags = 2.339244347e-06 wags = 7.881364039e-06 pags = -1.464004191e-11
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.800918564e-02 lketa = -1.410205681e-07 wketa = -7.128004331e-07 pketa = 1.212092823e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.669042343e-01 lpclm = 5.133079576e-08 wpclm = -3.307035300e-06 ppclm = 1.224487646e-12
+ pdiblc1 = 5.338088926e-01 lpdiblc1 = -2.875120856e-07 wpdiblc1 = -6.913575944e-07 ppdiblc1 = 1.382207041e-12
+ pdiblc2 = 2.028946854e-04 lpdiblc2 = 2.269383922e-10 wpdiblc2 = -1.019017709e-09 ppdiblc2 = 1.018268731e-15
+ pdiblcb = -6.114440459e-02 lpdiblcb = 1.191771629e-07 wpdiblcb = 4.173996457e-07 ppdiblcb = -8.345749362e-13
+ drout = -9.783071290e-02 ldrout = 1.315177920e-06 wdrout = 2.590144511e-06 pdrout = -5.178385265e-12
+ pscbe1 = 8.026643230e+08 lpscbe1 = -2.662364688e+00 wpscbe1 = -1.872036442e+01 ppscbe1 = 1.870660496e-5
+ pscbe2 = 6.541865313e-09 lpscbe2 = 2.295698733e-15 wpscbe2 = 1.193933210e-14 ppscbe2 = -1.007016969e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.533779899e-03 lalpha0 = 5.494187937e-09 walpha0 = 3.888206481e-08 palpha0 = -3.860387863e-14
+ alpha1 = 3.513156000e-10 walpha1 = -1.765821816e-15
+ beta0 = -8.141766918e+01 lbeta0 = 4.177076809e-05 wbeta0 = 6.126292737e-04 pbeta0 = -2.721582176e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.370713865e-10 lagidl = -3.704413905e-17 wagidl = -1.863323549e-16 pagidl = 1.861954006e-22
+ bgidl = -1.197910611e+08 lbgidl = 5.596663357e+02 wbgidl = 6.979565707e+03 pbgidl = -2.156171963e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.547960416e-01 lkt1 = -9.263619771e-08 wkt1 = -2.508082909e-07 pkt1 = 8.648669504e-14
+ kt2 = -1.145894977e-02 lkt2 = -3.725083360e-08 wkt2 = -2.019745422e-07 pkt2 = 2.127160445e-13
+ at = 1.316887331e+05 lat = 1.086190965e-01 wat = -6.763598968e-01 pat = 1.605292486e-8
+ ute = 5.199314551e-01 lute = -1.870448290e-06 wute = 3.910541676e-06 pute = -4.320061376e-12
+ ua1 = 2.941611603e-09 lua1 = -4.226664130e-15 wua1 = 9.639394328e-15 pua1 = -5.116115169e-21
+ ub1 = -1.751557943e-20 lub1 = 1.892396087e-24 wub1 = -1.418455486e-23 pub1 = 6.366960054e-30
+ uc1 = -6.972070325e-10 luc1 = 6.115133051e-16 wuc1 = 3.884635063e-15 puc1 = -3.284952573e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.14 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.075340383e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.985016835e-09 wvth0 = -1.638546819e-07 pvth0 = 1.914055131e-13
+ k1 = 4.363496353e-01 lk1 = 1.651807397e-08 wk1 = -1.862390226e-07 pk1 = 1.279476629e-13
+ k2 = 4.392349927e-02 lk2 = -1.427823290e-08 wk2 = -4.814891073e-08 pk2 = 2.594947727e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.736496513e+00 ldsub = -3.677069316e-07 wdsub = -5.174854288e-06 pdsub = 2.583623626e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.624903581e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.437367938e-08 wvoff = 2.544172144e-07 pvoff = -2.793379817e-13
+ nfactor = {-2.394520251e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.302947490e-06 wnfactor = 2.125508025e-05 pnfactor = -1.741821003e-11
+ eta0 = 5.260594773e-01 leta0 = -3.066019701e-07 weta0 = -7.095429572e-07 peta0 = 7.128788689e-13
+ etab = 1.521359777e+00 letab = -7.611588450e-07 wetab = -1.069657477e-05 petab = 5.348139527e-12
+ u0 = 1.260138607e-02 lu0 = 1.895392581e-10 wu0 = 7.530659612e-09 pu0 = -1.945918931e-14
+ ua = -1.592147237e-09 lua = 6.740884332e-16 wua = 7.464716430e-15 pua = -6.201309924e-21
+ ub = 2.854217280e-18 lub = -1.018814264e-24 wub = -9.324629433e-24 pub = 5.516381803e-30
+ uc = -1.390794640e-10 luc = 5.680197477e-17 wuc = 1.834588697e-16 puc = -5.504259020e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.082034147e+05 lvsat = -1.790097293e-01 wvsat = -1.281903781e+00 pvsat = 9.979269488e-7
+ a0 = 5.631264342e+00 la0 = -2.502465062e-06 wa0 = -2.316481008e-05 pa0 = 1.319636301e-11
+ ags = 3.354777145e+00 lags = -1.416006782e-06 wags = -1.645148853e-05 pags = 9.674926019e-12
+ a1 = 0.0
+ a2 = 1.769525333e-01 la2 = 6.225895268e-07 wa2 = 2.974599388e-06 pa2 = -2.972413057e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.990721982e-01 lketa = 8.589391091e-08 wketa = 1.025798870e-06 pketa = -5.252286103e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.992268668e-01 lpclm = 5.186644204e-07 wpclm = 3.926994178e-07 ppclm = -2.472527767e-12
+ pdiblc1 = 1.290551844e+00 lpdiblc1 = -1.043698831e-06 wpdiblc1 = -4.620926858e-06 ppdiblc1 = 5.308888072e-12
+ pdiblc2 = 2.165047594e-03 lpdiblc2 = -1.733772334e-09 wpdiblc2 = -1.462305453e-08 ppdiblc2 = 1.461230659e-14
+ pdiblcb = 1.411186489e-01 lpdiblcb = -8.293722725e-08 wpdiblcb = -8.349641585e-07 ppdiblcb = 4.168683806e-13
+ drout = 8.634212229e-01 ldrout = 3.546325046e-07 wdrout = -8.268904082e-07 pdrout = -1.763861867e-12
+ pscbe1 = 9.439485084e+08 lpscbe1 = -1.438427062e+02 wpscbe1 = -7.235301152e+02 ppscbe1 = 7.229983205e-4
+ pscbe2 = 8.938204582e-09 lpscbe2 = -9.887922620e-17 wpscbe2 = 9.476020178e-16 ppscbe2 = 9.134814632e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -7.104936726e-05 lalpha0 = 3.547251227e-11 walpha0 = 4.992157244e-10 palpha0 = -2.492409386e-16
+ alpha1 = 6.022617661e-10 lalpha1 = -2.507617206e-16 walpha1 = -3.529047874e-15 palpha1 = 1.761930087e-21
+ beta0 = -8.802961394e+01 lbeta0 = 4.837785308e-05 wbeta0 = 6.786283708e-04 pbeta0 = -3.381088054e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -2.987931674e+08 lbgidl = 7.385368754e+02 wbgidl = 9.716108970e+03 pbgidl = -4.890703868e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.070587498e-01 lkt1 = -4.041190260e-08 wkt1 = -3.116097251e-07 pkt1 = 1.472434402e-13
+ kt2 = -6.870796889e-02 lkt2 = 1.995610749e-08 wkt2 = 4.933925386e-08 pkt2 = -3.841303594e-14
+ at = 4.672041340e+05 lat = -2.266497006e-01 wat = -1.507385638e+00 pat = 8.464678619e-7
+ ute = -2.591959670e+00 lute = 1.239155594e-06 wute = -8.247878948e-07 pute = 4.117877283e-13
+ ua1 = -5.279442944e-09 lua1 = 3.988347942e-15 wua1 = 1.003213758e-14 pua1 = -5.508569758e-21
+ ub1 = 6.230931178e-18 lub1 = -4.351458062e-24 wub1 = -1.842492065e-23 pub1 = 1.060420918e-29
+ uc1 = 5.824814356e-11 luc1 = -1.433866114e-16 wuc1 = 9.577895785e-16 puc1 = -3.602583206e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.15 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.087849127e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.260161062e-09 wvth0 = 2.897461657e-07 pvth0 = -3.506151408e-14
+ k1 = 2.255219188e-01 lk1 = 1.217769739e-07 wk1 = -9.218370609e-08 pk1 = 8.098913524e-14
+ k2 = 9.826408992e-02 lk2 = -4.140858789e-08 wk2 = 6.074420956e-08 pk2 = -2.841704643e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.411559694e+00 ldsub = -2.054773508e-07 wdsub = -6.745863797e-07 pdsub = 3.367973689e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-9.274455099e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.037446100e-08 wvoff = -6.580303664e-07 pvoff = 1.762151597e-13
+ nfactor = {5.513335951e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.451683367e-07 wnfactor = -2.099604720e-05 pnfactor = 3.676299125e-12
+ eta0 = -6.643949407e-01 leta0 = 2.877502549e-07 weta0 = 1.434515617e-06 peta0 = -3.575745354e-13
+ etab = -5.765461730e-03 letab = 1.281337193e-09 wetab = 3.085650045e-08 petab = -7.691445584e-15
+ u0 = 2.103197838e-02 lu0 = -4.019560413e-09 wu0 = -6.354390936e-08 pu0 = 1.602585536e-14
+ ua = 1.558673532e-09 lua = -8.990060982e-16 wua = -1.101922003e-14 pua = 3.027072610e-21
+ ub = -2.489565998e-19 lub = 5.304918431e-25 wub = 4.462779592e-24 pub = -1.367188963e-30
+ uc = -8.456852788e-11 luc = 2.958657227e-17 wuc = 3.851451930e-16 puc = -1.557375124e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.981224373e+05 lvsat = 7.378104720e-02 wvsat = 1.538536824e+00 pvsat = -4.102203301e-7
+ a0 = 3.618937938e-01 la0 = 1.283472249e-07 wa0 = 7.188398290e-06 pa0 = -1.957931569e-12
+ ags = -2.123734998e+00 lags = 1.319222584e-06 wags = 1.188757757e-05 pags = -4.473777821e-12
+ a1 = 0.0
+ a2 = 2.046094933e+00 la2 = -3.106078536e-07 wa2 = -5.949198775e-06 pa2 = 1.482927033e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.814836225e-04 lketa = -1.398589053e-08 wketa = 1.744542395e-07 pketa = -1.001820333e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.140059907e+00 lpclm = -3.005460872e-07 wpclm = -7.619543551e-06 ppclm = 1.527704718e-12
+ pdiblc1 = -2.105346049e+00 lpdiblc1 = 6.517541305e-07 wpdiblc1 = 1.294985901e-05 ppdiblc1 = -3.463590333e-12
+ pdiblc2 = -1.090715258e-02 lpdiblc2 = 4.792719687e-09 wpdiblc2 = 2.819221161e-08 ppdiblc2 = -6.763857264e-15
+ pdiblcb = -0.025
+ drout = 2.286829735e+00 ldrout = -3.560255461e-07 wdrout = -6.630482921e-06 pdrout = 1.133668749e-12
+ pscbe1 = 5.121029832e+08 lpscbe1 = 7.176264989e+01 wpscbe1 = 1.447060230e+03 ppscbe1 = -3.607014683e-4
+ pscbe2 = 1.645755394e-08 lpscbe2 = -3.853027182e-15 wpscbe2 = 5.546343938e-15 ppscbe2 = -1.382509422e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.482740788e-08 lalpha0 = 2.742333230e-14 walpha0 = 2.760822894e-13 palpha0 = -1.378382242e-19
+ alpha1 = 4.502827321e-10 lalpha1 = -1.748839083e-16 walpha1 = -1.760630300e-15 palpha1 = 8.790210867e-22
+ beta0 = -1.851109849e+01 lbeta0 = 1.366969146e-05 wbeta0 = 1.406970190e-04 pbeta0 = -6.953850903e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.008731026e+09 lbgidl = 8.573580889e+01 wbgidl = 6.142080545e+02 pbgidl = -3.464433068e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.303376551e-01 lkt1 = -2.878955993e-08 wkt1 = -3.762461119e-07 pkt1 = 1.795141258e-13
+ kt2 = -2.366706548e-02 lkt2 = -2.531239153e-09 wkt2 = -2.324471784e-08 pkt2 = -2.174399301e-15
+ at = -3.869877714e+04 lat = 2.592991636e-02 wat = 5.159236304e-01 pat = -1.636996399e-7
+ ute = -1.121909516e-01 lute = 1.093865455e-09 wute = -4.049449690e-07 pute = 2.021748499e-13
+ ua1 = 4.278317483e-09 lua1 = -7.835073177e-16 wua1 = -2.475859766e-15 pua1 = 7.362355384e-22
+ ub1 = -4.588151770e-18 lub1 = 1.050131386e-24 wub1 = 8.196941801e-24 pub1 = -2.687154980e-30
+ uc1 = -3.290978658e-10 luc1 = 5.000169397e-17 wuc1 = 9.089174786e-17 puc1 = 7.255342478e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.16 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.907567519e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.194156981e-08 wvth0 = 6.867649150e-07 pvth0 = -1.340243926e-13
+ k1 = -5.534261136e-01 lk1 = 3.159414552e-07 wk1 = 4.875521954e-06 pk1 = -1.157286016e-12
+ k2 = 3.554480103e-01 lk2 = -1.055155378e-07 wk2 = -1.473253867e-06 pk2 = 3.539549841e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.443862747e+00 ldsub = -7.120593713e-07 wdsub = -1.726233469e-05 pdsub = 4.471542452e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.466105661e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.694754876e-08 wvoff = -1.657457231e-07 pvoff = 5.350582810e-14
+ nfactor = {8.911162818e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.492127651e-06 wnfactor = -4.745987326e-05 pnfactor = 1.027280473e-11
+ eta0 = 0.49
+ etab = -6.249997301e-04 letab = -6.727867937e-17 wetab = -1.356643062e-15 petab = 3.381636325e-22
+ u0 = 2.680577762e-02 lu0 = -5.458766479e-09 wu0 = -1.211807175e-07 pu0 = 3.039269435e-14
+ ua = 4.014747562e-09 lua = -1.511219391e-15 wua = -3.467453591e-14 pua = 8.923514924e-21
+ ub = -2.249249008e-18 lub = 1.029094730e-24 wub = 2.483811519e-23 pub = -6.446046990e-30
+ uc = 6.591225998e-11 luc = -7.923021318e-18 wuc = -2.657614586e-16 puc = 6.510734097e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.323662052e+05 lvsat = -3.352470427e-02 wvsat = -1.105344803e+00 pvsat = 2.488068237e-7
+ a0 = 3.464134057e+00 la0 = -6.449326942e-07 wa0 = -1.566094471e-05 pa0 = 3.737609913e-12
+ ags = 8.082407560e+00 lags = -1.224811541e-06 wags = -2.158029710e-05 pags = 3.868591960e-12
+ a1 = 0.0
+ a2 = -3.436580327e-03 la2 = 2.002686192e-07 wa2 = 7.002147203e-06 pa2 = -1.745390223e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.358819826e-01 lketa = -9.746486341e-08 wketa = -2.961905264e-06 pketa = 6.816026185e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.201693494e+00 lpclm = -6.664418348e-08 wpclm = -3.028023514e-06 ppclm = 3.831994765e-13
+ pdiblc1 = 8.820662159e-01 lpdiblc1 = -9.290318760e-08 wpdiblc1 = -4.153747715e-06 ppdiblc1 = 7.997401964e-13
+ pdiblc2 = 5.442631469e-03 lpdiblc2 = 7.172907656e-10 wpdiblc2 = 9.293908621e-09 ppdiblc2 = -2.053171769e-15
+ pdiblcb = 8.150898792e-01 lpdiblcb = -2.094050037e-07 wpdiblcb = -3.196628654e-06 ppdiblcb = 7.968076413e-13
+ drout = 4.968874310e-01 ldrout = 9.014442226e-08 wdrout = 4.590250026e-08 pdrout = -5.305204632e-13
+ pscbe1 = 7.986550012e+08 lpscbe1 = 3.352611287e-01 wpscbe1 = 1.129043578e+01 ppscbe1 = -2.814310474e-6
+ pscbe2 = -5.802180431e-08 lpscbe2 = 1.471207005e-14 wpscbe2 = 2.656766747e-13 ppscbe2 = -6.622389631e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.660659745e-08 lalpha0 = -2.845915044e-15 walpha0 = -3.342829089e-13 palpha0 = 1.430445694e-20
+ alpha1 = -2.513156000e-10 walpha1 = 1.765821816e-15
+ beta0 = 4.247839173e+01 lbeta0 = -1.532853821e-06 wbeta0 = -1.731330698e-04 pbeta0 = 8.688348043e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -9.644869147e+08 lbgidl = 5.775899789e+02 wbgidl = 1.271712259e+04 pbgidl = -3.363276298e-3
+ cgidl = 2.557872548e+03 lcgidl = -5.628086007e-04 wcgidl = -1.134877188e-02 pcgidl = 2.828851623e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.248335767e-01 lkt1 = -3.016153404e-08 wkt1 = -1.319410801e-07 pkt1 = 1.186174321e-13
+ kt2 = 1.551216517e-02 lkt2 = -1.229725008e-08 wkt2 = -1.138356271e-07 pkt2 = 2.040674369e-14
+ at = 1.158613815e+05 lat = -1.259652157e-02 wat = -2.752919108e-01 pat = 3.352270199e-8
+ ute = -1.480468140e+00 lute = 3.421574787e-07 wute = 1.215512015e-05 pute = -2.928609782e-12
+ ua1 = 3.074789045e-09 lua1 = -4.835098015e-16 wua1 = 1.701290771e-15 pua1 = -3.049818900e-22
+ ub1 = -1.516564861e-18 lub1 = 2.844922753e-25 wub1 = -9.199204028e-24 pub1 = 1.649095310e-30
+ uc1 = -4.336222390e-10 luc1 = 7.605596186e-17 wuc1 = 1.360136519e-15 puc1 = -2.438248730e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.17 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-7.460077387e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.205799066e-08 wvth0 = -1.730930487e-06 pvth0 = 3.277748379e-13
+ k1 = 2.116349876e+00 lk1 = -1.780808724e-07 wk1 = -1.177796127e-05 pk1 = 2.001462499e-12
+ k2 = -2.784739039e-02 lk2 = -4.029428105e-08 wk2 = 1.734361622e-06 pk2 = -2.420215262e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.339236393e+00 ldsub = 9.442297994e-07 wdsub = 5.144406113e-05 pdsub = -8.589074468e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.175493556e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.046271630e-09 wvoff = 1.651888621e-06 pvoff = -2.981581292e-13
+ nfactor = {-1.747570182e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.545189375e-06 wnfactor = 9.841734614e-05 pnfactor = -1.738360047e-11
+ eta0 = 1.985368093e+00 leta0 = -2.934884187e-07 weta0 = 7.145108178e-09 peta0 = -1.402334657e-15
+ etab = 3.254806901e-01 letab = -6.400313330e-08 wetab = -9.194629724e-07 petab = 1.804584004e-13
+ u0 = -7.031658291e-02 lu0 = 1.308528965e-08 wu0 = 4.595965323e-07 pu0 = -8.071136251e-14
+ ua = -2.545281267e-08 lua = 4.128919854e-15 wua = 1.440273573e-13 pua = -2.530318028e-20
+ ub = 2.038357293e-17 lub = -3.315345292e-24 wub = -1.120971704e-22 pub = 1.981826741e-29
+ uc = 2.911880464e-10 luc = -5.288812690e-17 wuc = -1.964386340e-15 puc = 3.405087703e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.071924122e+05 lvsat = 2.993956395e-02 wvsat = 2.049130203e+00 pvsat = -3.467114457e-7
+ a0 = -7.612516603e-01 la0 = 1.232025867e-07 wa0 = 1.006431457e-05 pa0 = -9.569142938e-13
+ ags = 1.25
+ a1 = 0.0
+ a2 = 3.034886182e+00 la2 = -3.770559894e-07 wa2 = -1.854008499e-05 pa2 = 3.102137703e-12
+ b0 = -4.103017639e-23 lb0 = 8.052787568e-30 wb0 = 2.062304679e-28 pb0 = -4.047582279e-35
+ b1 = 0.0
+ keta = -1.050643564e+00 lketa = 1.654188168e-07 wketa = 4.171961541e-06 pketa = -6.538882328e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.933750539e+00 lpclm = -2.166413389e-07 wpclm = -5.712175733e-06 ppclm = 9.463440595e-13
+ pdiblc1 = 1.010501991e+00 lpdiblc1 = -1.269207997e-07 wpdiblc1 = 4.680626576e-06 ppdiblc1 = -8.582975724e-13
+ pdiblc2 = 3.372419059e-02 lpdiblc2 = -4.765367551e-09 wpdiblc2 = 3.285536060e-08 ppdiblc2 = -6.872165858e-15
+ pdiblcb = -2.549616022e+00 lpdiblcb = 4.311107730e-07 wpdiblcb = 1.642347219e-05 ppdiblcb = -2.978368849e-12
+ drout = 9.983193450e-01 ldrout = 2.794341050e-10 wdrout = -1.906071842e-05 pdrout = 3.169130347e-12
+ pscbe1 = 8.034359437e+08 lpscbe1 = -5.712771792e-01 wpscbe1 = -2.884262897e+01 ppscbe1 = 4.795519705e-6
+ pscbe2 = 1.029119068e-07 lpscbe2 = -1.547841453e-14 wpscbe2 = -6.669319027e-13 ppscbe2 = 1.105344032e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.235866774e-07 lalpha0 = -3.392549333e-14 walpha0 = -1.123313769e-12 palpha0 = 1.705201142e-19
+ alpha1 = -2.513156000e-10 walpha1 = 1.765821816e-15
+ beta0 = 6.515295212e+01 lbeta0 = -6.128439510e-06 wbeta0 = -2.530473748e-04 pbeta0 = 2.519665970e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 4.768816516e+09 lbgidl = -4.928829945e+02 wbgidl = -1.928738887e+04 pbgidl = 2.599144022e-3
+ cgidl = -5.467977555e+03 lcgidl = 9.590127882e-04 wcgidl = 2.899165480e-02 pcgidl = -4.820297486e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.374254526e-01 lkt1 = 4.795554173e-08 wkt1 = 2.669070812e-06 pkt1 = -4.198744774e-13
+ kt2 = -8.082105042e-01 lkt2 = 1.482045108e-07 wkt2 = 4.818666436e-06 pkt2 = -9.457355680e-13
+ at = 4.354136266e+05 lat = -7.650799219e-02 wat = -2.506530004e+00 pat = 4.746156604e-7
+ ute = 5.303216873e+00 lute = -9.567950938e-07 wute = -3.403236030e-05 pute = 5.858651102e-12
+ ua1 = -2.949702508e-09 lua1 = 6.530349894e-16 wua1 = 2.200489760e-14 pua1 = -4.318791228e-21
+ ub1 = 4.975444341e-18 lub1 = -9.626830321e-25 wub1 = -3.010017501e-23 pub1 = 5.907610848e-30
+ uc1 = 5.118535911e-10 luc1 = -1.022953378e-16 wuc1 = -2.601343932e-15 puc1 = 5.105527668e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.18 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.108371908e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.416181897e-07 wvth0 = -1.804389422e-08 pvth0 = 1.804376160e-12
+ k1 = 4.567274430e-01 lk1 = -2.015547484e-06 wk1 = -9.830154391e-08 pk1 = 9.830082139e-12
+ k2 = 2.009262379e-02 lk2 = 8.988298148e-07 wk2 = 4.149548468e-08 pk2 = -4.149517969e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.324404127e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.153236349e-09 wvoff = 2.966567061e-09 pvoff = -2.966545257e-13
+ nfactor = {1.417739051e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.367127682e-06 wnfactor = -1.107518243e-07 pnfactor = 1.107510102e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.468976196e-02 lu0 = 2.446342401e-08 wu0 = 2.775832234e-09 pu0 = -2.775811832e-13
+ ua = -6.257063996e-10 lua = 5.242904420e-15 wua = 1.565995700e-16 pua = -1.565984190e-20
+ ub = 1.842195493e-18 lub = -3.894347687e-24 wub = 1.934507419e-25 pub = -1.934493201e-29
+ uc = -8.841333872e-11 luc = 1.074256376e-15 wuc = 5.636589784e-17 puc = -5.636548355e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.099215104e+05 lvsat = -9.921437448e-1
+ a0 = 1.413456932e+00 la0 = 6.435759524e-06 wa0 = 1.084107183e-07 pa0 = -1.084099215e-11
+ ags = 3.693493536e-01 lags = 4.480011712e-06 wags = 5.222966951e-08 pags = -5.222928563e-12
+ a1 = 0.0
+ a2 = 1.049985663e+00 la2 = -4.999529512e-6
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.193870672e-03 lketa = -1.636283240e-06 wketa = -3.585088859e-08 pketa = 3.585062509e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.877744279e-03 lpclm = 6.861141342e-06 wpclm = 2.192491956e-07 ppclm = -2.192475841e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 4.538491415e-03 lpdiblc2 = -9.108853203e-08 wpdiblc2 = -2.293044008e-10 ppdiblc2 = 2.293027154e-14
+ pdiblcb = 1.227248390e-03 lpdiblcb = -1.322982705e-07 wpdiblcb = -2.918457171e-09 ppdiblcb = 2.918435721e-13
+ drout = 0.56
+ pscbe1 = 7.804608126e+08 lpscbe1 = -3.398543280e+03 wpscbe1 = -1.359764284e+02 ppscbe1 = 1.359754290e-2
+ pscbe2 = 9.387568040e-09 lpscbe2 = 1.174235965e-14 wpscbe2 = 4.646520226e-16 ppscbe2 = -4.646486074e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.353153947e-10 lalpha0 = 2.353136651e-14 walpha0 = 7.121378026e-16 palpha0 = -7.121325684e-20
+ alpha1 = 1.626536487e-10 lalpha1 = -6.265318820e-15 walpha1 = -1.896094889e-16 palpha1 = 1.896080953e-20
+ beta0 = 5.105529510e+00 lbeta0 = -3.131381086e-05 wbeta0 = 4.083717435e-07 pbeta0 = -4.083687419e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.173748675e-10 lagidl = -1.737473978e-15 wagidl = -8.733150496e-17 pagidl = 8.733086307e-21
+ bgidl = 9.100775221e+08 lbgidl = 2.443652818e+04 wbgidl = 8.563761125e+02 pbgidl = -8.563698182e-2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.532117692e-01 lkt1 = 1.152168452e-06 wkt1 = 4.534668863e-08 pkt1 = -4.534635533e-12
+ kt2 = -0.037961
+ at = 0.0
+ ute = -2.801840520e-01 lute = -2.047579754e-06 wute = -4.000395509e-08 pute = 4.000366106e-12
+ ua1 = 2.320354091e-09 lua1 = -1.087532913e-14 wua1 = -5.466319908e-16 pua1 = 5.466279731e-20
+ ub1 = -1.049428527e-18 lub1 = 2.558366465e-23 wub1 = 1.445466103e-24 pub1 = -1.445455479e-28
+ uc1 = 2.356135282e-10 luc1 = -1.157626773e-14 wuc1 = -5.818636110e-16 puc1 = 5.818593343e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.19 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.115453077e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 7.217822942e-8
+ k1 = 3.559463651e-01 wk1 = 3.932206265e-7
+ k2 = 6.503576619e-02 wk2 = -1.659880388e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.322327432e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff = -1.186670435e-8
+ nfactor = {1.299378317e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 4.430235782e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.591297812e-02 wu0 = -1.110373700e-8
+ ua = -3.635515443e-10 wua = -6.264213011e-16
+ ub = 1.647470953e-18 wub = -7.738314060e-25
+ uc = -3.469854589e-11 wuc = -2.254718775e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.735256734e+00 wa0 = -4.336588101e-7
+ ags = 5.933581715e-01 wags = -2.089263561e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -7.862329813e-02 wketa = 1.434088246e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.499474192e-01 wpclm = -8.770290132e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.610256741e-05 wpdiblc2 = 9.172513120e-10
+ pdiblcb = -5.387908240e-03 wpdiblcb = 1.167425771e-8
+ drout = 0.56
+ pscbe1 = 6.105274035e+08 wpscbe1 = 5.439257030e+2
+ pscbe2 = 9.974707600e-09 wpscbe2 = -1.858676397e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.041296171e-09 walpha0 = -2.848655899e-15
+ alpha1 = -1.506238052e-10 walpha1 = 7.584658293e-16
+ beta0 = 3.539781426e+00 wbeta0 = -1.633547007e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.049797584e-11 wagidl = 3.493388580e-16
+ bgidl = 2.131948835e+09 wbgidl = -3.425630342e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.956012294e-01 wkt1 = -1.813934207e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.825668022e-01 wute = 1.600217011e-7
+ ua1 = 1.776567650e-09 wua1 = 2.186608321e-15
+ ub1 = 2.298017174e-19 wub1 = -5.782076905e-24
+ uc1 = -3.432211307e-10 wuc1 = 2.327539981e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.20 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.124951460e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.598007592e-08 wvth0 = 8.469359645e-08 pvth0 = -1.001137374e-13
+ k1 = 2.586802866e-01 lk1 = 7.780571373e-07 wk1 = 5.856805620e-07 pk1 = -1.539538026e-12
+ k2 = 1.029733714e-01 lk2 = -3.034729575e-07 wk2 = -2.429411810e-07 pk2 = 6.155685773e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.193889105e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.027412212e-07 wvoff = -4.934330307e-08 pvoff = 2.997852445e-13
+ nfactor = {1.580368183e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.247712400e-06 wnfactor = -6.637395005e-08 pnfactor = 4.074805819e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.502569979e-02 lu0 = 7.097574470e-09 wu0 = -2.946657669e-10 pu0 = -8.646462518e-14
+ ua = -7.404640344e-10 lua = 3.015022889e-15 wua = 1.965803097e-15 pua = -2.073588990e-20
+ ub = 1.955638623e-18 lub = -2.465114861e-24 wub = -2.003260352e-24 pub = 9.834527937e-30
+ uc = 4.610662326e-11 luc = -6.463819615e-16 wuc = -5.705315687e-16 puc = 2.760223911e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.308886950e+05 lvsat = -5.645576863e-01 wvsat = -2.866500015e-02 pvsat = 2.292989324e-7
+ a0 = 1.416770249e+00 la0 = 2.547657790e-06 wa0 = 7.114313066e-07 pa0 = -9.159879292e-12
+ ags = 3.594061272e-01 lags = 1.871444400e-06 wags = 4.215098314e-07 pags = -5.043026129e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.545708206e-02 lketa = -1.053200514e-07 wketa = 8.475269807e-08 pketa = 4.692059003e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.713431488e-02 lpclm = 2.262296967e-06 wpclm = -1.753896872e-06 ppclm = 7.014298375e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.471626697e-04 lpdiblc2 = 1.848310989e-09 wpdiblc2 = 1.834334079e-09 ppdiblc2 = -7.335988081e-15
+ pdiblcb = -7.069110030e-03 lpdiblcb = 1.344837864e-08 wpdiblcb = 2.005232279e-08 ppdiblcb = -6.701836275e-14
+ drout = 0.56
+ pscbe1 = 6.120625738e+08 lpscbe1 = -1.228023389e+01 wpscbe1 = 5.098077258e+02 ppscbe1 = 2.729187406e-4
+ pscbe2 = 1.167613135e-08 lpscbe2 = -1.361013948e-14 wpscbe2 = -7.637395898e-15 ppscbe2 = 4.622550865e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.982419379e-09 lalpha0 = -7.528293939e-15 walpha0 = -5.696788357e-15 palpha0 = 2.278296629e-20
+ alpha1 = -4.012015583e-10 lalpha1 = 2.004437850e-15 walpha1 = 1.516792290e-15 palpha1 = -6.066054319e-21
+ beta0 = 2.206423642e+00 lbeta0 = 1.066588225e-05 wbeta0 = -8.770178318e-06 pbeta0 = 5.708780506e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -9.447362404e-09 lagidl = 7.581591682e-14 wagidl = 2.917127997e-14 pagidl = -2.305543448e-19
+ bgidl = 9.830795530e+08 lbgidl = 9.190109835e+03 wbgidl = -5.487832968e+02 pbgidl = -2.301266188e-2
+ cgidl = 300.0
+ egidl = -4.271194736e-01 legidl = 4.216568356e-06 wegidl = 1.595227988e-06 pegidl = -1.276065141e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.028460191e-01 lkt1 = -7.419735073e-07 wkt1 = -6.277597631e-07 pkt1 = 3.570602659e-12
+ kt2 = -3.137221091e-02 lkt2 = -5.270546994e-8
+ at = -1.885734942e+05 lat = 1.508449352e+00 wat = 2.783135968e-02 pat = -2.226304214e-7
+ ute = 9.857563251e-01 lute = -1.094557930e-05 wute = -2.489888741e-06 pute = 2.119733586e-11
+ ua1 = 3.890536787e-09 lua1 = -1.691019933e-14 wua1 = 4.372814853e-15 pua1 = -1.748804539e-20
+ ub1 = -9.265925207e-20 lub1 = 2.579450747e-24 wub1 = -1.252433785e-23 pub1 = 5.393313199e-29
+ uc1 = -7.470080519e-10 luc1 = 3.229998586e-15 wuc1 = 4.654652277e-15 puc1 = -1.861518794e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.21 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.108119146e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.663192830e-09 wvth0 = 3.686263401e-08 pvth0 = 9.117495656e-14
+ k1 = 2.330764490e-01 lk1 = 8.804536689e-07 wk1 = 1.104870565e-06 pk1 = -3.615916433e-12
+ k2 = 1.073118101e-01 lk2 = -3.208235234e-07 wk2 = -4.182256280e-07 pk2 = 1.316577531e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.475001779e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.683186368e-09 wvoff = 6.034968894e-10 pvoff = 1.000347556e-13
+ nfactor = {1.086688735e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.733574615e-07 wnfactor = 4.707496751e-07 pnfactor = 1.926706104e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.583991471e-02 lu0 = -3.615133676e-08 wu0 = -5.372633934e-08 pu0 = 1.272227968e-13
+ ua = 1.780324383e-09 lua = -7.066278002e-15 wua = -1.001031237e-14 pua = 2.715976953e-20
+ ub = 6.325522522e-19 lub = 2.826258155e-24 wub = 3.733125986e-24 pub = -1.310680117e-29
+ uc = -2.090406046e-10 luc = 3.740194168e-16 wuc = 4.301543582e-16 puc = -1.241784292e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.707457297e+05 lvsat = -3.240300302e-01 wvsat = -7.809866016e-02 pvsat = 4.269972387e-7
+ a0 = 1.741258866e+00 la0 = 1.249941821e-06 wa0 = 5.120339004e-07 pa0 = -8.362436224e-12
+ ags = -2.794610997e-02 lags = 3.420568645e-06 wags = 2.366073129e-06 pags = -1.281985007e-11
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.672382567e-02 lketa = -2.202319580e-07 wketa = -1.375005123e-08 pketa = 8.631444980e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.182328751e-01 lpclm = 5.830778362e-08 wpclm = 9.592234190e-07 ppclm = -3.836188647e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -4.135226813e-02 lpdiblcb = 1.505558129e-07 wpdiblcb = 1.849336478e-07 ppdiblcb = -7.264224752e-13
+ drout = 0.56
+ pscbe1 = 4.193862592e+08 lpscbe1 = 7.582834076e+02 wpscbe1 = 1.151855931e+03 ppscbe1 = -2.294802176e-3
+ pscbe2 = -2.628972864e-09 lpscbe2 = 4.359976314e-14 wpscbe2 = 5.866591313e-14 ppscbe2 = -2.189389945e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.784652266e-03 lalpha0 = 1.113656275e-08 walpha0 = 8.427226872e-09 palpha0 = -3.370271348e-14
+ alpha1 = 3.512232415e-10 lalpha1 = -1.004708317e-15 walpha1 = -7.602799105e-16 palpha1 = 3.040560836e-21
+ beta0 = -6.452983849e+01 lbeta0 = 2.775618796e-04 wbeta0 = 2.121139034e-04 pbeta0 = -8.262861719e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.891674225e-08 lagidl = -3.761965420e-14 wagidl = -5.694533289e-14 pagidl = 1.138488110e-19
+ bgidl = 5.105698789e+09 lbgidl = -7.297336982e+03 wbgidl = -1.199319565e+04 pbgidl = 2.275657589e-2
+ cgidl = 300.0
+ egidl = 1.154238947e+00 legidl = -2.107703029e-06 wegidl = -3.190455977e-06 pegidl = 6.378566969e-12
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.584975230e-01 lkt1 = 2.804446043e-07 wkt1 = 6.516046036e-07 pkt1 = -1.545914474e-12
+ kt2 = -3.976450213e-02 lkt2 = -1.914247339e-08 wkt2 = -1.168823923e-09 pkt2 = 4.674436607e-15
+ at = 3.704577405e+05 lat = -7.272646985e-01 wat = -2.885977421e-01 pat = 1.042853410e-6
+ ute = -3.332000681e+00 lute = 6.322275174e-06 wute = 5.106426196e-06 pute = -9.182340603e-12
+ ua1 = -2.337184545e-09 lua1 = 7.996108623e-15 wua1 = -2.883185176e-15 pua1 = 1.153062156e-20
+ ub1 = 2.085743962e-18 lub1 = -6.132560983e-24 wub1 = 3.318139585e-24 pub1 = -9.425133521e-30
+ uc1 = 2.779738022e-11 luc1 = 1.313463398e-16 wuc1 = 1.952935112e-16 puc1 = -7.810305039e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.22 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.120937485e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.429045049e-08 wvth0 = 1.005694963e-07 pvth0 = -3.619194346e-14
+ k1 = 9.180689596e-01 lk1 = -4.890278829e-07 wk1 = -1.470372633e-06 pk1 = 1.532677159e-12
+ k2 = -1.366451056e-01 lk2 = 1.669109996e-07 wk2 = 5.063842648e-07 pk2 = -5.319626662e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.066573261e-02 ldsub = 9.583162241e-07 wdsub = 9.358283226e-07 pdsub = -1.870968811e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.701779398e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.502204201e-08 wvoff = 1.412592791e-07 pvoff = -1.811734268e-13
+ nfactor = {2.749730633e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.349477270e-06 wnfactor = 2.635705169e-06 pnfactor = -2.401613642e-12
+ eta0 = -6.141591779e-02 leta0 = 2.827278949e-07 weta0 = 7.634052067e-09 peta0 = -1.526249311e-14
+ etab = -6.365577510e-01 letab = 1.132699082e-06 wetab = 4.021299398e-06 petab = -8.039643142e-12
+ u0 = 3.645452315e-03 lu0 = 8.221275094e-09 wu0 = 2.713145092e-08 pu0 = -3.443335320e-14
+ ua = -3.151877288e-09 lua = 2.794500172e-15 wua = 8.712505697e-15 pua = -1.027210534e-20
+ ub = 3.237495007e-18 lub = -2.381712722e-24 wub = -6.767194413e-24 pub = 7.886121892e-30
+ uc = 2.547668733e-11 luc = -9.484279684e-17 wuc = -4.457844803e-16 puc = 5.094495696e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.449722111e+04 lvsat = 1.462829678e-01 wvsat = 3.169817455e-01 pvsat = -3.628731885e-7
+ a0 = 3.547777757e+00 la0 = -2.361768168e-06 wa0 = -7.144693865e-06 pa0 = 6.945391612e-12
+ ags = 2.803491073e+00 lags = -2.240224616e-06 wags = -8.236647350e-06 pags = 8.377797892e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.821275787e-01 lketa = 2.703951763e-07 wketa = 8.460437073e-07 pketa = -8.558110707e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.188999078e-01 lpclm = -1.429522914e-07 wpclm = -2.060488178e-06 ppclm = 2.201015059e-12
+ pdiblc1 = 3.769820107e-01 lpdiblc1 = 2.602641031e-08 wpdiblc1 = 9.690324363e-08 ppdiblc1 = -1.937352634e-13
+ pdiblc2 = 1.580250000e-07 lpdiblc2 = 4.295260411e-10
+ pdiblcb = 9.286329557e-02 lpdiblcb = -1.177766660e-07 wpdiblcb = -3.566911057e-07 ppdiblcb = 3.564289378e-13
+ drout = 8.525995111e-01 ldrout = -5.849839615e-07 wdrout = -2.187014329e-06 pdrout = 4.372421203e-12
+ pscbe1 = 7.973356770e+08 lpscbe1 = 2.662364688e+00 wpscbe1 = 8.063072563e+00 ppscbe1 = -8.057146204e-6
+ pscbe2 = 2.925890079e-08 lpscbe2 = -2.015254659e-14 wpscbe2 = -1.022435759e-13 ppscbe2 = 1.027617152e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.533780099e-03 lalpha0 = -5.494187937e-09 walpha0 = -1.674694482e-08 palpha0 = 1.662712689e-14
+ alpha1 = -1.513156000e-10 walpha1 = 7.605594161e-16
+ beta0 = 9.143480343e+01 lbeta0 = -3.425277020e-05 wbeta0 = -2.561811836e-04 pbeta0 = 1.099598052e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.268158399e+09 lbgidl = 3.749232047e+02 wbgidl = 3.298679380e+00 pbgidl = -1.227595347e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.447457429e-01 lkt1 = -1.469018482e-07 wkt1 = -3.013242275e-07 pkt1 = 3.592427852e-13
+ kt2 = -3.819969981e-02 lkt2 = -2.227092790e-08 wkt2 = -6.756718940e-08 pkt2 = 1.374223648e-13
+ at = -1.051779731e+05 lat = 2.236571364e-01 wat = 5.142060712e-01 pat = -5.621641555e-7
+ ute = 3.261939694e+00 lute = -6.860759031e-06 wute = -9.871647240e-06 pute = 2.076279739e-11
+ ua1 = 7.935435959e-09 lua1 = -1.254158201e-14 wua1 = -1.546112496e-14 pua1 = 3.667725634e-20
+ ub1 = -4.824276575e-18 lub1 = 7.682401227e-24 wub1 = 9.975725618e-24 pub1 = -2.273541226e-29
+ uc1 = -4.312723030e-11 luc1 = 2.731434313e-16 wuc1 = 5.970259038e-16 puc1 = -1.584200016e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.23 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.133869556e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.721301581e-08 wvth0 = 1.303312005e-07 pvth0 = -6.593177279e-14
+ k1 = 5.035933658e-01 lk1 = -7.485692862e-08 wk1 = -5.242269920e-07 pk1 = 5.872269349e-13
+ k2 = -7.467799960e-03 lk2 = 3.782863928e-08 wk2 = 2.101597933e-07 pk2 = -2.359559197e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.079315335e+00 ldsub = -3.959937062e-08 wdsub = -1.871656645e-06 pdsub = 9.344526549e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.913819039e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.371607880e-08 wvoff = -1.029960624e-07 pvoff = 6.290238693e-14
+ nfactor = {2.468084280e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.420220100e-07 wnfactor = -3.185887255e-06 pnfactor = 3.415699912e-12
+ eta0 = 4.207248234e-01 leta0 = -1.990584729e-07 weta0 = -1.800981224e-07 peta0 = 1.723316982e-13
+ etab = 9.927769337e-01 letab = -4.954380417e-07 wetab = -8.039752481e-06 petab = 4.012543864e-12
+ u0 = 1.861199518e-02 lu0 = -6.734267367e-09 wu0 = -2.268053711e-08 pu0 = 1.534202301e-14
+ ua = 5.761459899e-10 lua = -9.307830084e-16 wua = -3.433801835e-15 pua = 1.865274661e-21
+ ub = 8.943319870e-19 lub = -4.027192674e-26 wub = 5.263655348e-25 pub = 5.979227107e-31
+ uc = -1.601071847e-10 luc = 9.060467105e-17 wuc = 2.891507548e-16 puc = -2.249454882e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.950388989e+04 lvsat = 1.238034763e-02 wvsat = -8.212549537e-02 pvsat = 3.594070856e-8
+ a0 = 9.662028680e-01 la0 = 2.179092630e-07 wa0 = 2.832443853e-07 pa0 = -4.770871040e-13
+ ags = 2.527917188e-01 lags = 3.085999748e-07 wags = -8.599419616e-07 pags = 1.006514383e-12
+ a1 = 0.0
+ a2 = 1.023655437e+00 la2 = -2.234910506e-07 wa2 = -1.281193579e-06 pa2 = 1.280251902e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.308885863e-02 lketa = 1.554199703e-09 wketa = 9.098857884e-08 pketa = -1.013109078e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.398163810e-01 lpclm = -6.392689108e-08 wpclm = -3.139473443e-07 ppclm = 4.557579327e-13
+ pdiblc1 = 1.321938900e+00 lpdiblc1 = -9.182359354e-07 wpdiblc1 = -4.778687995e-06 ppdiblc1 = 4.678272415e-12
+ pdiblc2 = -1.633322462e-03 lpdiblc2 = 2.061805920e-09 wpdiblc2 = 4.468738464e-09 ppdiblc2 = -4.465453942e-15
+ pdiblcb = 1.226899351e-02 lpdiblcb = -3.724160080e-08 wpdiblcb = -1.873255893e-07 ppdiblcb = 1.871879050e-13
+ drout = 2.289163275e-01 ldrout = 3.824081491e-08 wdrout = 2.362329162e-06 pdrout = -1.735785205e-13
+ pscbe1 = 7.867858752e+08 lpscbe1 = 1.320441242e+01 wpscbe1 = 6.641831408e+01 ppscbe1 = -6.636949662e-5
+ pscbe2 = 8.807320979e-09 lpscbe2 = 2.840013135e-16 wpscbe2 = 1.605463840e-15 ppscbe2 = -1.010995588e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.104956726e-05 lalpha0 = -3.547251227e-11 walpha0 = -2.150178554e-10 palpha0 = 1.073508896e-16
+ alpha1 = -4.022617661e-10 lalpha1 = 2.507617206e-16 walpha1 = 1.520000810e-15 palpha1 = -7.588832043e-22
+ beta0 = 1.052920706e+02 lbeta0 = -4.809985232e-05 wbeta0 = -2.930667322e-04 pbeta0 = 1.468182430e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 2.168329474e+09 lbgidl = -5.245862443e+02 wbgidl = -2.684419167e+03 pbgidl = 1.458147026e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.923368963e-01 lkt1 = 5.808256884e-10 wkt1 = 1.170248461e-07 pkt1 = -5.879880189e-14
+ kt2 = -1.069128953e-01 lkt2 = 4.639176342e-08 wkt2 = 2.413691341e-07 pkt2 = -1.712868906e-13
+ at = 1.628938226e+05 lat = -4.421762657e-02 wat = 2.217293220e-02 pat = -7.049266085e-8
+ ute = -6.956611576e+00 lute = 3.350281604e-06 wute = 2.111331436e-05 pute = -1.019939027e-11
+ ua1 = -1.227173678e-08 lua1 = 7.650738462e-15 wua1 = 4.517758801e-14 pua1 = -2.391688718e-20
+ ub1 = 8.024857567e-18 lub1 = -5.157288802e-24 wub1 = -2.744175438e-23 pub1 = 1.465456589e-29
+ uc1 = 8.105819158e-10 luc1 = -5.799382386e-16 wuc1 = -2.823674689e-15 puc1 = 1.833986362e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.24 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.022957729e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.161377518e-09 wvth0 = -3.641824747e-08 pvth0 = 1.732039034e-14
+ k1 = -1.800998899e-01 lk1 = 2.664871847e-07 wk1 = 1.946598058e-06 pk1 = -6.463695338e-13
+ k2 = 2.546118198e-01 lk2 = -9.301854207e-08 wk2 = -7.251082612e-07 pk2 = 2.309906856e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.072479709e+00 ldsub = -3.618658192e-08 wdsub = 1.029735420e-06 pdsub = -5.141108545e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.160152022e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.141753511e-08 wvoff = -3.843361293e-08 pvoff = 3.066861562e-14
+ nfactor = {1.036183838e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.271242354e-07 wnfactor = 1.507516187e-06 pnfactor = 1.072447842e-12
+ eta0 = -4.445805757e-01 leta0 = 2.329582272e-07 weta0 = 3.296600365e-07 peta0 = -8.217270900e-14
+ etab = 1.506098876e-03 letab = -5.312083614e-10 wetab = -5.692631887e-09 petab = 1.418973887e-15
+ u0 = 7.760312850e-03 lu0 = -1.316402186e-09 wu0 = 3.163622373e-09 pu0 = 2.438938728e-15
+ ua = 8.482032857e-11 lua = -6.854813021e-16 wua = -3.611173982e-15 pua = 1.953830365e-21
+ ub = -6.256339584e-19 lub = 7.185938710e-25 wub = 6.356077519e-24 pub = -2.312648443e-30
+ uc = 4.716850742e-11 luc = -1.288082738e-17 wuc = -2.770062483e-16 puc = 5.771688802e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.372788543e+04 lvsat = 2.861544911e-04 wvsat = 7.160604496e-02 pvsat = -4.081206893e-8
+ a0 = 2.106991064e+00 la0 = -3.516463557e-07 wa0 = -1.583005060e-06 pa0 = 4.546659255e-13
+ ags = 2.335674504e-01 lags = 3.181979791e-07 wags = 3.903998637e-08 pags = 5.576841604e-13
+ a1 = 0.0
+ a2 = 3.526891253e-01 la2 = 1.114989452e-07 wa2 = 2.562387159e-06 pa2 = -6.387134352e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.301051841e-01 lketa = -6.993757402e-08 wketa = -4.745617655e-07 pketa = 1.810485849e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.874294788e-01 lpclm = 6.208105566e-08 wpclm = 1.189723801e-06 ppclm = -2.949724415e-13
+ pdiblc1 = -1.268767243e+00 lpdiblc1 = 3.752129670e-07 wpdiblc1 = 8.744952916e-06 ppdiblc1 = -2.073608164e-12
+ pdiblc2 = -4.295785301e-03 lpdiblc2 = 3.391080429e-09 wpdiblc2 = -5.038583098e-09 ppdiblc2 = 2.812189581e-16
+ pdiblcb = -9.953798701e-02 lpdiblcb = 1.857971133e-08 wpdiblcb = 3.746511786e-07 ppdiblcb = -9.338742603e-14
+ drout = 1.584293583e-01 ldrout = 7.343249158e-08 wdrout = 4.067521432e-06 pdrout = -1.024921339e-12
+ pscbe1 = 8.262059567e+08 lpscbe1 = -6.476654557e+00 wpscbe1 = -1.317193145e+02 ppscbe1 = 3.255368652e-5
+ pscbe2 = 3.000980360e-08 lpscbe2 = -1.030165617e-14 wpscbe2 = -6.257149115e-14 ppscbe2 = 3.103031185e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.929962619e+00 lbeta0 = 1.037554125e-08 wbeta0 = 2.769684253e-06 pbeta0 = -8.825255295e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 7.979420898e+08 lbgidl = 1.596002130e+02 wbgidl = 1.673699015e+03 pbgidl = -7.177088475e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.222934637e-01 lkt1 = 1.553709128e-08 wkt1 = 8.595247211e-08 pkt1 = -4.328545307e-14
+ kt2 = -2.548854002e-03 lkt2 = -5.713549675e-09 wkt2 = -1.293914376e-07 pkt2 = 1.382088627e-14
+ at = 1.211319864e+05 lat = -2.336740344e-02 wat = -2.874356545e-01 pat = 8.408407019e-8
+ ute = -4.239885812e-01 lute = 8.877158429e-08 wute = 1.162247198e-06 pute = -2.385207203e-13
+ ua1 = 5.699153929e-09 lua1 = -1.321498289e-15 wua1 = -9.617427042e-15 pua1 = 3.440346014e-21
+ ub1 = -4.553389348e-18 lub1 = 1.122589644e-24 wub1 = 8.022215023e-24 pub1 = -3.051352793e-30
+ uc1 = -7.464764405e-10 luc1 = 1.974465016e-16 wuc1 = 2.188766686e-15 puc1 = -6.685501814e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.25 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.430731570e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.300030531e-08 wvth0 = -5.553891022e-08 pvth0 = 2.208650234e-14
+ k1 = 1.133504781e+00 lk1 = -6.094848361e-08 wk1 = -3.603519045e-06 pk1 = 7.370804060e-13
+ k2 = -1.650048527e-01 lk2 = 1.157720780e-08 wk2 = 1.142704604e-06 pk2 = -2.345896882e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -9.549673461e-01 ldsub = 4.691850083e-07 wdsub = 4.847557791e-06 pdsub = -1.465760348e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.586452320e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.913607461e-10 wvoff = 3.973754625e-07 pvoff = -7.796333357e-14
+ nfactor = {-4.780393732e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.322744973e-06 wnfactor = 2.135816173e-05 pnfactor = -3.875623318e-12
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = -1.239046954e-02 lu0 = 3.706482586e-09 wu0 = 7.583184992e-08 pu0 = -1.567470701e-14
+ ua = -7.549987824e-09 lua = 1.217609152e-15 wua = 2.345343234e-14 pua = -4.792428728e-21
+ ub = 6.160584680e-18 lub = -9.729729178e-25 wub = -1.743233280e-23 pub = 3.616969654e-30
+ uc = 1.057282890e-10 luc = -2.747773134e-17 wuc = -4.658892432e-16 puc = 1.047988078e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.610851531e+04 lvsat = 4.678046784e-03 wvsat = -3.199449009e-01 pvsat = 5.678787761e-8
+ a0 = -3.675973068e-01 la0 = 2.651819146e-07 wa0 = 3.598532628e-06 pa0 = -8.369100663e-13
+ ags = 2.176241710e+00 lags = -1.660427201e-07 wags = 8.105935181e-06 pags = -1.453110470e-12
+ a1 = 0.0
+ a2 = 1.750539365e+00 la2 = -2.369361948e-07 wa2 = -1.813883138e-06 pa2 = 4.521375804e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.574068287e-01 lketa = 1.014351078e-07 wketa = 1.528043007e-06 pketa = -3.181306938e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.121649329e-01 lpclm = -6.871712730e-08 wpclm = -1.572762631e-06 ppclm = 3.936187389e-13
+ pdiblc1 = -1.045740275e-01 lpdiblc1 = 8.502034512e-08 wpdiblc1 = 8.054139805e-07 ppdiblc1 = -9.455899122e-14
+ pdiblc2 = 1.341439983e-02 lpdiblc2 = -1.023448866e-09 wpdiblc2 = -3.077468633e-08 ppdiblc2 = 6.696328731e-15
+ pdiblcb = -2.855674619e-01 lpdiblcb = 6.495034839e-08 wpdiblcb = 2.335618548e-06 ppdiblcb = -5.821879573e-13
+ drout = 1.561647109e+00 ldrout = -2.763405809e-07 wdrout = -5.305911845e-06 pdrout = 1.311547506e-12
+ pscbe1 = 8.030589294e+08 lpscbe1 = -7.069108033e-01 wpscbe1 = -1.084508145e+01 ppscbe1 = 2.423970813e-6
+ pscbe2 = -2.611671098e-08 lpscbe2 = 3.688719486e-15 wpscbe2 = 1.053117212e-13 ppscbe2 = -1.081709708e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.887686193e+00 lbeta0 = 2.701785748e-07 wbeta0 = 7.306085555e-07 pbeta0 = -3.742553258e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 9.546499493e-10 lagidl = -2.130343196e-16 wagidl = -4.295737296e-15 pagidl = 1.070776957e-21
+ bgidl = 2.206765983e+09 lbgidl = -1.915702746e+02 wbgidl = -3.222583903e+03 pbgidl = 5.027631141e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.981906457e-01 lkt1 = 9.529102359e-09 wkt1 = 2.367744361e-07 pkt1 = -8.088008993e-14
+ kt2 = 6.189064144e-02 lkt2 = -2.177606051e-08 wkt2 = -3.469483189e-07 pkt2 = 6.805020229e-14
+ at = -4.461763687e+04 lat = 1.794817641e-02 wat = 5.313257048e-01 pat = -1.200044800e-7
+ ute = 2.279410999e+00 lute = -5.850913121e-07 wute = -6.743205482e-06 pute = 1.732031942e-12
+ ua1 = 2.292349755e-09 lua1 = -4.723012466e-16 wua1 = 5.634074764e-15 pua1 = -3.613195839e-22
+ ub1 = -2.448570693e-18 lub1 = 5.979320224e-25 wub1 = -4.514651931e-24 pub1 = 7.364934814e-32
+ uc1 = 1.209712750e-10 luc1 = -1.877785315e-17 wuc1 = -1.427423516e-15 puc1 = 2.328394693e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.26 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-1.088774217e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.803894332e-09 wvth0 = -8.079221129e-09 pvth0 = 1.486632645e-14
+ k1 = -9.839013862e-01 lk1 = 3.488443911e-07 wk1 = 3.804868851e-06 pk1 = -6.470282759e-13
+ k2 = 5.532753209e-01 lk2 = -1.282981645e-07 wk2 = -1.186542436e-06 pk2 = 2.003134492e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 9.184455469e+00 ldsub = -1.476335211e-06 wdsub = -2.155654556e-05 pdsub = 3.577440490e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.800711661e-03+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.088346659e-08 wvoff = 7.489004668e-08 pvoff = -2.206412685e-14
+ nfactor = {3.407135859e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.587424030e-07 wnfactor = -6.546311486e-06 pnfactor = 1.233516271e-12
+ eta0 = 1.987245422e+00 leta0 = -2.938568727e-07 weta0 = -2.290932418e-09 peta0 = 4.496298511e-16
+ etab = 3.607201594e-01 letab = -7.091940770e-08 wetab = -1.096587539e-06 petab = 2.152217534e-13
+ u0 = 3.556478130e-02 lu0 = -5.353962771e-09 wu0 = -7.259623919e-08 pu0 = 1.197007320e-14
+ ua = 7.449175569e-09 lua = -1.610733737e-15 wua = -2.134830106e-14 pua = 3.546109438e-21
+ ub = -5.244867779e-18 lub = 1.173249559e-24 wub = 1.671936871e-23 pub = -2.742810756e-30
+ uc = -2.502241278e-10 luc = 3.977751048e-17 wuc = 7.569201675e-16 puc = -1.252576349e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.878749816e+05 lvsat = -3.644067172e-02 wvsat = 6.339822036e-02 pvsat = -1.306367061e-8
+ a0 = 3.164905054e+00 la0 = -4.029770165e-07 wa0 = -9.669774041e-06 pa0 = 1.687828560e-12
+ ags = 1.25
+ a1 = 0.0
+ a2 = -1.822583639e+00 la2 = 4.418737356e-07 wa2 = 5.875073854e-06 pa2 = -1.014058600e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.951101457e-02 lketa = -1.395031161e-08 wketa = -1.508547977e-06 pketa = 2.476769696e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.661291027e-03 lpclm = 1.032700448e-07 wpclm = 3.994081330e-06 ppclm = -6.616303672e-13
+ pdiblc1 = 1.654926791e+00 lpdiblc1 = -2.522454613e-07 wpdiblc1 = 1.441546471e-06 ppdiblc1 = -2.283767220e-13
+ pdiblc2 = 3.275687064e-02 lpdiblc2 = -4.916754269e-09 wpdiblc2 = 3.771741247e-08 ppdiblc2 = -6.111248979e-15
+ pdiblcb = -5.524661761e+00 lpdiblcb = 1.099360541e-06 wpdiblcb = 3.137698029e-05 ppdiblcb = -6.337200678e-12
+ drout = -5.410491700e+00 ldrout = 1.065840402e-06 wdrout = 1.315196544e-05 pdrout = -2.186711535e-12
+ pscbe1 = 7.942137480e+08 lpscbe1 = 9.620511823e-01 wpscbe1 = 1.751100374e+01 ppscbe1 = -2.911467038e-6
+ pscbe2 = -8.910157842e-08 lpscbe2 = 1.640025194e-14 wpscbe2 = 2.981877823e-13 ppscbe2 = -4.969772063e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.607287247e+01 lbeta0 = -1.310665523e-06 wbeta0 = -6.355581455e-06 pbeta0 = 9.810244976e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.823217985e-09 lagidl = 3.119615294e-16 wagidl = 9.666693636e-15 pagidl = -1.568015979e-21
+ bgidl = 8.279294079e+08 lbgidl = 6.088015590e+01 wbgidl = 5.207392976e+02 pbgidl = -1.842423464e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.781271391e-01 lkt1 = -5.238450104e-08 wkt1 = -6.447682126e-07 pkt1 = 8.446588371e-14
+ kt2 = 4.155326256e-01 lkt2 = -9.324866480e-08 wkt2 = -1.332248343e-06 pkt2 = 2.678834261e-13
+ at = -7.996610376e+04 lat = 2.658789887e-02 wat = 8.392931885e-02 pat = -4.357645405e-8
+ ute = -5.830121880e+00 lute = 9.510409699e-07 wute = 2.192727387e-05 pute = -3.730728199e-12
+ ua1 = -1.353329944e-09 lua1 = 1.984289618e-16 wua1 = 1.398103103e-14 pua1 = -2.033799496e-21
+ ub1 = 9.095071142e-19 lub1 = -4.438224060e-27 wub1 = -9.663505934e-24 pub1 = 1.091173470e-30
+ uc1 = 2.601997860e-11 luc1 = -1.922972210e-18 wuc1 = -1.593926157e-16 puc1 = 6.049941308e-24
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.27 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.136357815e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.950664129e-07 wvth0 = 6.665019407e-08 pvth0 = -1.332954893e-12
+ k1 = 4.303063649e-01 lk1 = 1.111437855e-06 wk1 = -1.834311824e-08 pk1 = 3.668488826e-13
+ k2 = 2.638046037e-02 lk2 = -3.238477856e-07 wk2 = 2.246652937e-08 pk2 = -4.493140746e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.259010590e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.050496832e-07 wvoff = -1.682355728e-08 pvoff = 3.364587804e-13
+ nfactor = {1.397729005e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.607625912e-07 wnfactor = -5.019518244e-08 pnfactor = 1.003866755e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.872379925e-02 lu0 = -1.295929703e-07 wu0 = -9.432423216e-09 pu0 = 1.886415315e-13
+ ua = -7.895001713e-10 lua = 4.378978693e-15 wua = 6.522906270e-16 pua = -1.304533311e-20
+ ub = 2.690642107e-18 lub = -2.597649106e-23 wub = -2.374213426e-24 pub = 4.748252348e-29
+ uc = -6.501065391e-11 luc = -8.838022409e-16 wuc = -1.445792803e-17 puc = 2.891479340e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.104448434e+05 lvsat = -3.002536521e+00 wvsat = -3.042149690e-01 pvsat = 6.084075782e-6
+ a0 = 1.015743251e+00 la0 = 1.152392345e-05 wa0 = 1.312016402e-06 pa0 = -2.623936371e-11
+ ags = 3.797879703e-02 lags = 9.726497598e-06 wags = 1.055060361e-06 pags = -2.110043176e-11
+ a1 = 0.0
+ a2 = 1.556534611e+00 la2 = -1.513013616e-05 wa2 = -1.532975160e-06 pa2 = 3.065837646e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = 8.486766206e-02 lketa = -2.321987405e-06 wketa = -2.830212636e-07 pketa = 5.660217251e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.738862078e-01 lpclm = 4.680475441e-06 wpclm = 7.662973128e-07 ppclm = -1.532538303e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.322952610e-02 lpdiblc2 = -2.588412182e-07 wpdiblc2 = -2.653108695e-08 ppdiblc2 = 5.306022387e-13
+ pdiblcb = 7.784338305e-03 lpdiblcb = -1.862863718e-07 wpdiblcb = -2.276225707e-08 ppdiblcb = 4.552284111e-13
+ drout = 0.56
+ pscbe1 = 8.057711559e+08 lpscbe1 = -3.102197179e+02 wpscbe1 = -2.125734242e+02 ppscbe1 = 4.251312243e-3
+ pscbe2 = 9.288006224e-09 lpscbe2 = 1.450532220e-15 wpscbe2 = 7.659571439e-16 ppscbe2 = -1.531857990e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.486805178e-10 lalpha0 = 1.897291308e-14 walpha0 = 2.871003235e-15 palpha0 = -5.741795451e-20
+ alpha1 = 3.525899165e-10 lalpha1 = -5.051612677e-15 walpha1 = -7.644158954e-16 palpha1 = 1.528775606e-20
+ beta0 = 9.236345025e+00 lbeta0 = -1.247223168e-04 wbeta0 = -1.209276482e-05 pbeta0 = 2.418464082e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.851746450e-11 lagidl = 1.148245110e-15
+ bgidl = 4.434138120e+08 lbgidl = 1.113131467e+04 wbgidl = 2.268646099e+03 pbgidl = -4.537125452e-2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.635563411e-01 lkt1 = 1.603209296e-07 wkt1 = 7.665259062e-08 pkt1 = -1.532995473e-12
+ kt2 = -0.037961
+ at = 0.0
+ ute = -1.665818966e-01 lute = -3.262042184e-06 wute = -3.837995212e-07 pute = 7.675708332e-12
+ ua1 = 2.139727641e-09 lua1 = 7.187183033e-15
+ ub1 = -2.501969717e-19 lub1 = -2.861100907e-23 wub1 = -9.732579431e-25 pub1 = 1.946444352e-29
+ uc1 = 4.334531165e-11 luc1 = 7.650412604e-15 puc1 = -3.308722450e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.28 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.09160285+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4858803
+ k2 = 0.010187476
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.23615392+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4457689+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0122439126
+ ua = -5.7054319e-10
+ ub = 1.39176982e-18
+ uc = -1.0920239e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.5919606
+ ags = 0.52432155
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.031235975
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.060146165
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 790259600.0
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.4593183e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.45554
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.29 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.096965714e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.289897344e-8
+ k1 = 4.522097581e-01 lk1 = 2.693395874e-7
+ k2 = 2.269705454e-02 lk2 = -1.000674338e-07 wk2 = 1.387778781e-23 pk2 = -5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.356936746e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.681625035e-9
+ nfactor = {1.558435894e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.012531388e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.492833185e-02 lu0 = -2.147338093e-8
+ ua = -9.089350183e-11 lua = -3.836844963e-15
+ ub = 1.293690895e-18 lub = 7.845593095e-25
+ uc = -1.424170877e-10 luc = 2.656931686e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.214167700e+05 lvsat = -4.887892486e-01 wvsat = -2.328306437e-16
+ a0 = 1.651852193e+00 la0 = -4.790887229e-7
+ ags = 4.986878111e-01 lags = 2.050510707e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.745180763e-02 lketa = 4.972209241e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.124149426e-01 lpclm = 4.580068028e-06 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 3.589658719e-04 lpdiblc2 = -5.757576728e-10
+ pdiblcb = -4.431168108e-04 lpdiblcb = -8.696847218e-9
+ drout = 0.56
+ pscbe1 = 7.805209898e+08 lpscbe1 = 7.790172373e+1
+ pscbe2 = 9.152466940e-09 lpscbe2 = 1.664395553e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -6.915519527e-01 lbeta0 = 2.952970233e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.918552200e-10 lagidl = -3.673533665e-16
+ bgidl = 8.017422366e+08 lbgidl = 1.585916388e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.102799397e-01 lkt1 = 4.378792836e-7
+ kt2 = -3.137221091e-02 lkt2 = -5.270546994e-8
+ at = -1.793770334e+05 lat = 1.434884425e+0
+ ute = 1.630094498e-01 lute = -3.941233465e-6
+ ua1 = 5.335468721e-09 lua1 = -2.268886504e-14
+ ub1 = -4.231141289e-18 lub1 = 2.040085581e-23
+ uc1 = 7.910528872e-10 luc1 = -2.921114695e-15 wuc1 = 8.271806126e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.30 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.095938434e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.879060751e-8
+ k1 = 5.981645711e-01 lk1 = -3.143723879e-7
+ k2 = -3.088465745e-02 lk2 = 1.142200316e-07 wk2 = 1.040834086e-23 pk2 = -2.081668171e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.473007613e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.273819047e-8
+ nfactor = {1.242240996e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.632940483e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.086841217e-03 lu0 = 5.887553094e-9
+ ua = -1.527435151e-09 lua = 1.908265777e-15
+ ub = 1.866108470e-18 lub = -1.504690264e-24
+ uc = -6.690246480e-11 luc = -3.630981963e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.449391836e+05 lvsat = -1.829351138e-1
+ a0 = 1.910452889e+00 la0 = -1.513301435e-6
+ ags = 7.538877290e-01 lags = -8.155610292e-07 wags = 8.881784197e-22
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.126732654e-02 lketa = 6.498136366e-08 wketa = 5.551115123e-23
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.351940539e-01 lpclm = -1.209303965e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = 1.975631812e-02 lpdiblcb = -8.947974034e-08 ppdiblcb = 4.163336342e-29
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.675630966e-08 lpscbe2 = -2.874538651e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.560060825e+00 lbeta0 = 4.527846154e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.142724829e+09 lbgidl = 2.222366395e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.431844278e-01 lkt1 = -2.303799486e-7
+ kt2 = -4.015072270e-02 lkt2 = -1.759787501e-8
+ at = 2.750948889e+05 lat = -3.826692271e-1
+ ute = -1.644657739e+00 lute = 3.288106654e-6
+ ua1 = -3.289890404e-09 lua1 = 1.180623182e-14 wua1 = 8.271806126e-31 pua1 = 4.963083675e-36
+ ub1 = 3.182174067e-18 lub1 = -9.246956829e-24 pub1 = -3.081487911e-45
+ uc1 = 9.232922993e-11 luc1 = -1.267336281e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.31 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.087705784e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.233135855e-8
+ k1 = 4.322060899e-01 lk1 = 1.742259510e-8
+ k2 = 3.068207834e-02 lk2 = -8.868188432e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.898963481e-01 ldsub = 3.400822775e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.235009021e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.844034868e-9
+ nfactor = {1.145902819e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.558995947e-7
+ eta0 = -5.889335829e-02 leta0 = 2.776846300e-7
+ etab = 6.922211054e-01 letab = -1.523881978e-06 wetab = 4.440892099e-22 petab = 1.110223025e-28
+ u0 = 1.261063863e-02 lu0 = -3.156716733e-9
+ ua = -2.729587568e-10 lua = -5.997649717e-16
+ ub = 1.001375792e-18 lub = 2.241395141e-25
+ uc = -1.218261949e-10 luc = 7.349727172e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.024470420e+04 lvsat = 2.637689452e-2
+ a0 = 1.186919436e+00 la0 = -6.676632695e-8
+ ags = 8.181288894e-02 lags = 5.280946760e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.564960161e-03 lketa = -1.239492287e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.804209211e-02 lpclm = 5.843405517e-7
+ pdiblc1 = 4.090022531e-01 lpdiblc1 = -3.799053949e-8
+ pdiblc2 = 1.580250000e-07 lpdiblc2 = 4.295260411e-10
+ pdiblcb = -0.025
+ drout = 1.299330017e-01 ldrout = 8.598178973e-7
+ pscbe1 = 800000000.0
+ pscbe2 = -4.525975301e-09 lpscbe2 = 1.380354094e-14 ppscbe2 = -6.617444900e-36
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.783523713e+00 lbeta0 = 2.081819624e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.269248399e+09 lbgidl = -3.071750489e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443138732e-01 lkt1 = -2.819538791e-8
+ kt2 = -6.052627731e-02 lkt2 = 2.313825818e-8
+ at = 6.473381100e+04 lat = 3.789831325e-2
+ ute = 0.0
+ ua1 = 2.826536098e-09 lua1 = -4.221256071e-16
+ ub1 = -1.527945722e-18 lub1 = 1.698208119e-25
+ uc1 = 1.541511415e-10 luc1 = -2.503320121e-16 wuc1 = 1.033975766e-31 puc1 = 1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.32 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.090803540e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.542683752e-8
+ k1 = 3.303703168e-01 lk1 = 1.191835189e-7
+ k2 = 6.197639260e-02 lk2 = -4.013950137e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.608541037e-01 ldsub = 2.691766759e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.254154280e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.930916229e-9
+ nfactor = {1.415355000e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.866454611e-7
+ eta0 = 3.612140650e-01 leta0 = -1.421140143e-7
+ etab = -1.663840256e+00 letab = 8.304476780e-7
+ u0 = 1.111754745e-02 lu0 = -1.664722981e-09 wu0 = -1.387778781e-23
+ ua = -5.585029939e-10 lua = -3.144306096e-16
+ ub = 1.068261686e-18 lub = 1.573027816e-25
+ uc = -6.456159825e-11 luc = 1.627476450e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.236673570e+04 lvsat = 2.425642272e-2
+ a0 = 1.059796782e+00 la0 = 6.026289207e-8
+ ags = -3.136337212e-02 lags = 6.411877525e-7
+ a1 = 0.0
+ a2 = 6.003039853e-01 la2 = 1.995492381e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.697697029e-02 lketa = -3.192249000e-08 pketa = -1.387778781e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.360771286e-01 lpclm = 8.667157091e-8
+ pdiblc1 = -2.571078061e-01 lpdiblc1 = 6.276299288e-7
+ pdiblc2 = -1.566939902e-04 lpdiblc2 = 5.862627701e-10
+ pdiblcb = -4.962997438e-02 lpdiblcb = 2.461187135e-8
+ drout = 1.009513028e+00 ldrout = -1.911563762e-8
+ pscbe1 = 8.087328239e+08 lpscbe1 = -8.726405225e+0
+ pscbe2 = 9.337822739e-09 lpscbe2 = -5.006721217e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.452507416e+00 lbeta0 = 4.140626236e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.281302899e+09 lbgidl = -4.276314530e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.536677683e-01 lkt1 = -1.884836796e-8
+ kt2 = -2.715603810e-02 lkt2 = -1.020745390e-8
+ at = 1.702205398e+05 lat = -6.751088280e-2
+ ute = 1.997060000e-02 lute = -1.995592161e-8
+ ua1 = 2.656528384e-09 lua1 = -2.522428491e-16
+ ub1 = -1.042863932e-18 lub1 = -3.149044430e-25
+ uc1 = -1.224595845e-10 luc1 = 2.607540497e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.33 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.034991600e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.438110935e-9
+ k1 = 4.631246217e-01 lk1 = 5.290394085e-8
+ k2 = 1.501052909e-02 lk2 = -1.669108952e-08 pk2 = -6.938893904e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.412740535e+00 ldsub = -2.060669031e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.287150206e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.283545090e-9
+ nfactor = {1.534320245e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.272502780e-7
+ eta0 = -3.356492968e-01 leta0 = 2.058054720e-07 weta0 = -2.220446049e-22 peta0 = 1.110223025e-28
+ etab = -3.749470590e-04 letab = -6.232944635e-11
+ u0 = 8.805685030e-03 lu0 = -5.104909885e-10
+ ua = -1.108438655e-09 lua = -3.986698167e-17
+ ub = 1.474637765e-18 lub = -4.558657148e-26
+ uc = -4.436410663e-11 luc = 6.190863850e-18 wuc = 5.169878828e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.173890430e+05 lvsat = -1.319958952e-2
+ a0 = 1.583910476e+00 la0 = -2.014087313e-7
+ ags = 2.464676360e-01 lags = 5.024764542e-7
+ a1 = 0.0
+ a2 = 1.199392029e+00 la2 = -9.955445421e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.670672610e-02 lketa = -1.011274932e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.805560965e-01 lpclm = -3.538822096e-8
+ pdiblc1 = 1.620872991e+00 lpdiblc1 = -3.099801539e-7
+ pdiblc2 = -5.960710496e-03 lpdiblc2 = 3.484005071e-09 ppdiblc2 = -8.673617380e-31
+ pdiblcb = 2.425994875e-02 lpdiblcb = -1.227878113e-08 wpdiblcb = 1.387778781e-23 ppdiblcb = -6.505213035e-31
+ drout = 1.502481601e+00 ldrout = -2.652375925e-7
+ pscbe1 = 7.826812591e+08 lpscbe1 = 4.280229240e+0
+ pscbe2 = 9.333980631e-09 lpscbe2 = -4.814898237e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.845163779e+00 lbeta0 = -2.812419554e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.350991152e+09 lbgidl = -7.755605097e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.938917417e-01 lkt1 = 1.234054096e-9
+ kt2 = -4.530433909e-02 lkt2 = -1.146642408e-9
+ at = 2.615312949e+04 lat = 4.416932803e-3
+ ute = -3.994120000e-02 lute = 9.955943218e-9
+ ua1 = 2.521217536e-09 lua1 = -1.846868784e-16
+ ub1 = -1.902567152e-18 lub1 = 1.143152850e-25
+ uc1 = -2.323089072e-11 luc1 = -2.346600883e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.34 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.614251969e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.570214029e-08 wvth0 = 8.839817767e-14 pvth0 = -2.203457239e-20
+ k1 = -5.722461056e-02 lk1 = 1.826087922e-07 wk1 = -3.987795658e-13 pk1 = 9.940178813e-20
+ k2 = 2.125849839e-01 lk2 = -6.593948599e-08 wk2 = -4.975484957e-14 pk2 = 1.240214262e-20
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.468363388e-01 ldsub = -1.515379369e-08 wdsub = 7.790399614e-14 pdsub = -1.941873995e-20
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.273383794e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.655319356e-08 wvoff = -4.098910811e-14 pvoff = 1.021715001e-20
+ nfactor = {2.277094436e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.210266923e-08 wnfactor = 5.931075009e-13 pnfactor = -1.478409430e-19
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 1.266704449e-02 lu0 = -1.472992754e-09 wu0 = -5.481675669e-15 pu0 = 1.366389887e-21
+ ua = 1.998517754e-10 lua = -3.659779959e-16 wua = -2.419839623e-22 pua = 6.031813269e-29
+ ub = 4.003284706e-19 lub = 2.222011347e-25 wub = -3.088505014e-31 pub = 7.698562060e-38
+ uc = -4.821791451e-11 luc = 7.151483271e-18 wuc = -7.407702238e-26 puc = 1.846480385e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.961254947e+04 lvsat = 2.344276242e-02 wvsat = 2.605019556e-08 pvsat = -6.493401946e-15
+ a0 = 8.214845247e-01 la0 = -1.136262656e-08 wa0 = 1.160535135e-14 pa0 = -2.892808659e-21
+ ags = 4.854727851e+00 lags = -6.462015284e-07 wags = 4.284101749e-13 pags = -1.067876632e-19
+ a1 = 0.0
+ a2 = 1.151168225e+00 la2 = -8.753394759e-08 wa2 = 9.353417774e-13 pa2 = -2.331479680e-19
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.248763730e-02 lketa = -3.686470494e-09 wketa = -6.173064282e-16 pketa = 1.538728589e-22
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.924688054e-01 lpclm = 6.134835765e-08 wpclm = -4.074220072e-15 ppclm = 1.015560525e-21
+ pdiblc1 = 1.615631159e-01 lpdiblc1 = 5.377472217e-08 wpdiblc1 = -5.000176806e-14 ppdiblc1 = 1.246369097e-20
+ pdiblc2 = 3.245360502e-03 lpdiblc2 = 1.189253784e-09 wpdiblc2 = -6.000212827e-16 ppdiblc2 = 1.495643123e-22
+ pdiblcb = 4.862030192e-01 lpdiblcb = -1.274250206e-07 wpdiblcb = 2.797629930e-13 ppdiblcb = -6.973512250e-20
+ drout = -1.916129469e-01 ldrout = 1.570408851e-07 wdrout = 1.004973864e-13 pdrout = -2.505048080e-20
+ pscbe1 = 7.994753355e+08 lpscbe1 = 9.405379727e-02 wpscbe1 = -8.148437500e-06 ppscbe1 = 2.031120300e-12
+ pscbe2 = 8.681988012e-09 lpscbe2 = 1.143699577e-16 wpscbe2 = 8.358320747e-22 ppscbe2 = -2.083436816e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.129104825e+00 lbeta0 = 1.465114798e-07 wbeta0 = 4.506332800e-13 pbeta0 = -1.123271005e-19
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.648127901e-10 lagidl = 1.407880601e-16 wagidl = -1.740802484e-22 pagidl = 4.339211319e-29
+ bgidl = 1.141910710e+09 lbgidl = -2.543961448e+01 wbgidl = 3.864334412e-04 pbgidl = -9.632433176e-11
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.199520018e-01 lkt1 = -1.719653517e-08 wkt1 = -1.108681200e-13 pkt1 = 2.763554185e-20
+ kt2 = -5.275329183e-02 lkt2 = 7.101207958e-10 wkt2 = -7.944725544e-15 pkt2 = 1.980342001e-21
+ at = 1.309510566e+05 lat = -2.170552250e-02 wat = 6.086635450e-08 pat = -1.517185185e-14
+ ute = 5.121857576e-02 lute = -1.276699829e-08 wute = -1.311157638e-14 pute = 3.268257068e-21
+ ua1 = 4.154046646e-09 lua1 = -5.916940266e-16 wua1 = -8.778088769e-22 pua1 = 2.188070291e-28
+ ub1 = -3.940370848e-18 lub1 = 6.222684232e-25 wub1 = 7.778053586e-31 pub1 = -1.938796520e-37
+ uc1 = -3.506996717e-10 luc1 = 5.816049688e-17 wuc1 = -6.975555789e-23 puc1 = 1.738761922e-29
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.35 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-1.091444326e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.891446422e-09 wvth0 = 1.359594393e-12 pvth0 = -2.736154725e-19
+ k1 = 2.733610754e-01 lk1 = 1.350434900e-07 wk1 = 3.765382743e-13 pk1 = -4.333952841e-20
+ k2 = 1.611999296e-01 lk2 = -6.210755014e-08 wk2 = 2.620938844e-14 pk2 = -1.330862531e-21
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.061414258e+00 ldsub = -2.942229886e-07 wdsub = -4.687326438e-13 pdsub = 8.602538859e-20
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {2.094558561e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.817422975e-08 wvoff = 3.028874573e-14 pvoff = -2.803288712e-21
+ nfactor = {1.244004252e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.488547807e-07 wnfactor = -3.455916016e-13 pnfactor = 2.237283425e-20
+ eta0 = 1.986488332e+00 leta0 = -2.937082825e-07 weta0 = 2.570175290e-13 peta0 = -5.044354578e-20
+ etab = -1.630959850e-03 letab = 1.974347099e-10 wetab = 8.810806217e-16 petab = -1.729252878e-22
+ u0 = 1.157642340e-02 lu0 = -1.398628374e-09 wu0 = 1.617483419e-14 pu0 = -2.754447982e-21
+ ua = 3.949451567e-10 lua = -4.389743043e-16 wua = 1.091251803e-21 pua = -1.956293183e-28
+ ub = 2.797998630e-19 lub = 2.669283874e-25 wub = 7.319085622e-31 pub = -1.199782819e-37
+ uc = -1.110656404e-13 luc = -1.612020295e-18 wuc = 6.313561129e-24 puc = -1.233453944e-30
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.088240009e+05 lvsat = -4.075737074e-02 wvsat = -4.810017860e-08 pvsat = 7.443940965e-15
+ a0 = -3.032888734e-02 la0 = 1.547409959e-07 wa0 = 7.787949912e-13 pa0 = -1.537396130e-19
+ ags = 1.250000362e+00 lags = -6.012721077e-14 wags = -1.094419730e-12 pags = 1.819636974e-19
+ a1 = 0.0
+ a2 = 1.187482526e-01 la2 = 1.067929675e-07 wa2 = -2.144329503e-12 pa2 = 3.491739031e-19
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.189664782e-01 lketa = 6.789090505e-08 wketa = 4.409042553e-13 pketa = -8.648676447e-20
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.322446062e+00 lpclm = -1.153558612e-07 wpclm = 8.403277079e-13 ppclm = -1.646146774e-19
+ pdiblc1 = 2.131264901e+00 lpdiblc1 = -3.277092517e-07 wpdiblc1 = -1.267594815e-12 ppdiblc1 = 2.526165424e-19
+ pdiblc2 = 4.522001127e-02 lpdiblc2 = -6.936122122e-09 wpdiblc2 = 6.042993089e-14 ppdiblc2 = -1.181429582e-20
+ pdiblcb = 4.843401116e+00 lpdiblcb = -9.946744331e-07 wpdiblcb = -1.281277469e-11 ppdiblcb = 2.493258689e-18
+ drout = -1.064619979e+00 ldrout = 3.432740603e-07 wdrout = 1.706933869e-12 pdrout = -3.427133155e-19
+ pscbe1 = 7.999999931e+08 lpscbe1 = 1.143630028e-06 wpscbe1 = 2.081605911e-05 ppscbe1 = -3.460982323e-12
+ pscbe2 = 9.430160657e-09 lpscbe2 = -2.162425182e-17 wpscbe2 = -2.068863309e-21 ppscbe2 = 3.419887848e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.397276455e+01 lbeta0 = -9.865004674e-07 wbeta0 = 3.351150895e-13 pbeta0 = -1.003070906e-19
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.370998103e-09 lagidl = -2.061661974e-16 wagidl = -8.404522904e-22 pagidl = 1.782925689e-28
+ bgidl = 1.000000326e+09 lbgidl = -5.423579121e-05 wbgidl = -9.871856689e-04 pbgidl = 1.641344252e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.911813583e-01 lkt1 = -2.447398172e-08 wkt1 = 3.278208176e-13 pkt1 = -5.584301777e-20
+ kt2 = -2.468915302e-02 lkt2 = -4.730545465e-09 wkt2 = 1.084893364e-13 pkt2 = -2.068379001e-20
+ at = -5.223289612e+04 lat = 1.218870496e-02 wat = -2.020222822e-08 pat = -6.996985612e-16
+ ute = 1.415421327e+00 lute = -2.817229670e-07 wute = -4.838224307e-13 pute = 9.596225700e-20
+ ua1 = 3.266493694e-09 lua1 = -4.736097814e-16 wua1 = 3.311341522e-21 pua1 = -5.826267374e-28
+ ub1 = -2.283654412e-18 lub1 = 3.561237281e-25 wub1 = -2.889616718e-30 pub1 = 5.075210096e-37
+ uc1 = -2.664901037e-11 luc1 = 7.615108932e-20 wuc1 = 1.776628973e-22 puc1 = -2.952306690e-29
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.36 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.103465450e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.372432872e-7
+ k1 = 4.212539000e-01 lk1 = 1.292480499e-6
+ k2 = 3.746785924e-02 lk2 = -5.455876137e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.342036093e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.900477982e-8
+ nfactor = {1.372957310e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.456178280e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.406882844e-02 lu0 = -3.649697542e-8
+ ua = -4.675899092e-10 lua = -2.058989945e-15
+ ub = 1.518950173e-18 lub = -2.543513577e-24 wub = 3.081487911e-39
+ uc = -7.214574862e-11 luc = -7.411055910e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.663233076e+00 la0 = -1.425397138e-6
+ ags = 5.586589101e-01 lags = -6.867219644e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.480543051e-02 lketa = 4.713717867e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.042871993e-01 lpclm = -2.882714742e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.362379205e-04 lpdiblc2 = 3.014921787e-9
+ pdiblcb = -3.449004373e-03 lpdiblcb = 3.837222522e-8
+ drout = 0.56
+ pscbe1 = 7.008645946e+08 lpscbe1 = 1.787834404e+3
+ pscbe2 = 9.666011755e-09 lpscbe2 = -6.109300570e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.681808713e-10 lalpha0 = -9.363273314e-15
+ alpha1 = -2.465499712e-11 lalpha1 = 2.493008321e-15 walpha1 = 1.050131637e-32 palpha1 = 5.557619741e-37
+ beta0 = 3.268475902e+00 lbeta0 = -5.369320704e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.851746450e-11 lagidl = 1.148245110e-15
+ bgidl = 1.563007487e+09 lbgidl = -1.125973593e+4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.257277191e-01 lkt1 = -5.962237055e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.559898067e-01 lute = 5.259768035e-7
+ ua1 = 2.139727641e-09 lua1 = 7.187183033e-15
+ ub1 = -7.305069847e-19 lub1 = -1.900516184e-23
+ uc1 = 4.334531165e-11 luc1 = 7.650412604e-15 puc1 = 6.617444900e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.37 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.09160285+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4858803
+ k2 = 0.010187476
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.23615392+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4457689+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0122439126
+ ua = -5.7054319e-10
+ ub = 1.39176982e-18
+ uc = -1.0920239e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.5919606
+ ags = 0.52432155
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.031235975
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.060146165
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 790259600.0
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.4593183e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.45554
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.38 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.096965714e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.289897344e-8
+ k1 = 4.522097581e-01 lk1 = 2.693395874e-7
+ k2 = 2.269705454e-02 lk2 = -1.000674338e-07 pk2 = -1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.356936746e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.681625035e-9
+ nfactor = {1.558435894e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.012531388e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.492833185e-02 lu0 = -2.147338093e-8
+ ua = -9.089350183e-11 lua = -3.836844963e-15
+ ub = 1.293690895e-18 lub = 7.845593095e-25
+ uc = -1.424170877e-10 luc = 2.656931686e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.214167700e+05 lvsat = -4.887892486e-1
+ a0 = 1.651852193e+00 la0 = -4.790887229e-7
+ ags = 4.986878111e-01 lags = 2.050510707e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.745180763e-02 lketa = 4.972209241e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.124149426e-01 lpclm = 4.580068028e-06 wpclm = 2.220446049e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.589658719e-04 lpdiblc2 = -5.757576728e-10
+ pdiblcb = -4.431168108e-04 lpdiblcb = -8.696847218e-9
+ drout = 0.56
+ pscbe1 = 7.805209898e+08 lpscbe1 = 7.790172373e+1
+ pscbe2 = 9.152466940e-09 lpscbe2 = 1.664395553e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -6.915519527e-01 lbeta0 = 2.952970233e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.918552200e-10 lagidl = -3.673533665e-16
+ bgidl = 8.017422366e+08 lbgidl = 1.585916388e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.102799397e-01 lkt1 = 4.378792836e-7
+ kt2 = -3.137221091e-02 lkt2 = -5.270546994e-8
+ at = -1.793770334e+05 lat = 1.434884425e+0
+ ute = 1.630094498e-01 lute = -3.941233465e-6
+ ua1 = 5.335468721e-09 lua1 = -2.268886504e-14 pua1 = 2.646977960e-35
+ ub1 = -4.231141289e-18 lub1 = 2.040085581e-23
+ uc1 = 7.910528872e-10 luc1 = -2.921114695e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.39 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.095938434e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.879060751e-8
+ k1 = 5.981645711e-01 lk1 = -3.143723879e-7
+ k2 = -3.088465745e-02 lk2 = 1.142200316e-07 wk2 = -1.387778781e-23 pk2 = -2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.473007613e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.273819047e-8
+ nfactor = {1.242240996e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.632940483e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.086841217e-03 lu0 = 5.887553094e-9
+ ua = -1.527435151e-09 lua = 1.908265777e-15
+ ub = 1.866108470e-18 lub = -1.504690264e-24
+ uc = -6.690246480e-11 luc = -3.630981963e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.449391836e+05 lvsat = -1.829351138e-1
+ a0 = 1.910452889e+00 la0 = -1.513301435e-6
+ ags = 7.538877290e-01 lags = -8.155610292e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.126732654e-02 lketa = 6.498136366e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.351940539e-01 lpclm = -1.209303965e-06 wpclm = 1.776356839e-21
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = 1.975631812e-02 lpdiblcb = -8.947974034e-08 wpdiblcb = -1.387778781e-23 ppdiblcb = -1.387778781e-29
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.675630966e-08 lpscbe2 = -2.874538651e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.560060825e+00 lbeta0 = 4.527846154e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.142724829e+09 lbgidl = 2.222366395e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.431844278e-01 lkt1 = -2.303799486e-7
+ kt2 = -4.015072270e-02 lkt2 = -1.759787501e-8
+ at = 2.750948889e+05 lat = -3.826692271e-1
+ ute = -1.644657739e+00 lute = 3.288106654e-6
+ ua1 = -3.289890404e-09 lua1 = 1.180623182e-14 pua1 = 1.654361225e-36
+ ub1 = 3.182174067e-18 lub1 = -9.246956829e-24 wub1 = -3.081487911e-39
+ uc1 = 9.232922993e-11 luc1 = -1.267336281e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.40 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.087705784e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.233135855e-8
+ k1 = 4.322060899e-01 lk1 = 1.742259510e-8
+ k2 = 3.068207834e-02 lk2 = -8.868188432e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.898963481e-01 ldsub = 3.400822775e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.235009021e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.844034868e-9
+ nfactor = {1.145902819e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.558995947e-7
+ eta0 = -5.889335829e-02 leta0 = 2.776846300e-07 peta0 = -2.220446049e-28
+ etab = 6.922211054e-01 letab = -1.523881978e-06 petab = 1.332267630e-27
+ u0 = 1.261063863e-02 lu0 = -3.156716733e-9
+ ua = -2.729587568e-10 lua = -5.997649717e-16
+ ub = 1.001375792e-18 lub = 2.241395141e-25
+ uc = -1.218261949e-10 luc = 7.349727172e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.024470420e+04 lvsat = 2.637689452e-2
+ a0 = 1.186919436e+00 la0 = -6.676632695e-8
+ ags = 8.181288894e-02 lags = 5.280946760e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.564960160e-03 lketa = -1.239492287e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.804209211e-02 lpclm = 5.843405517e-7
+ pdiblc1 = 4.090022531e-01 lpdiblc1 = -3.799053949e-8
+ pdiblc2 = 1.580250000e-07 lpdiblc2 = 4.295260411e-10
+ pdiblcb = -0.025
+ drout = 1.299330017e-01 ldrout = 8.598178973e-7
+ pscbe1 = 800000000.0
+ pscbe2 = -4.525975301e-09 lpscbe2 = 1.380354094e-14 ppscbe2 = 6.617444900e-36
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.783523713e+00 lbeta0 = 2.081819624e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.269248399e+09 lbgidl = -3.071750489e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443138732e-01 lkt1 = -2.819538791e-8
+ kt2 = -6.052627731e-02 lkt2 = 2.313825818e-8
+ at = 6.473381100e+04 lat = 3.789831325e-2
+ ute = 0.0
+ ua1 = 2.826536098e-09 lua1 = -4.221256071e-16 wua1 = -6.617444900e-30
+ ub1 = -1.527945722e-18 lub1 = 1.698208119e-25
+ uc1 = 1.541511415e-10 luc1 = -2.503320121e-16 wuc1 = 1.033975766e-31 puc1 = -2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.41 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.090803540e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.542683752e-8
+ k1 = 3.303703168e-01 lk1 = 1.191835189e-7
+ k2 = 6.197639260e-02 lk2 = -4.013950137e-08 wk2 = 5.551115123e-23 pk2 = 2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.608541037e-01 ldsub = 2.691766759e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.254154280e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.930916229e-9
+ nfactor = {1.415355000e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.866454611e-7
+ eta0 = 3.612140650e-01 leta0 = -1.421140143e-7
+ etab = -1.663840256e+00 letab = 8.304476780e-7
+ u0 = 1.111754745e-02 lu0 = -1.664722981e-9
+ ua = -5.585029939e-10 lua = -3.144306096e-16
+ ub = 1.068261686e-18 lub = 1.573027816e-25
+ uc = -6.456159825e-11 luc = 1.627476450e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.236673570e+04 lvsat = 2.425642272e-2
+ a0 = 1.059796782e+00 la0 = 6.026289207e-8
+ ags = -3.136337212e-02 lags = 6.411877525e-7
+ a1 = 0.0
+ a2 = 6.003039853e-01 la2 = 1.995492381e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.697697029e-02 lketa = -3.192249000e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.360771286e-01 lpclm = 8.667157091e-8
+ pdiblc1 = -2.571078061e-01 lpdiblc1 = 6.276299288e-7
+ pdiblc2 = -1.566939902e-04 lpdiblc2 = 5.862627701e-10
+ pdiblcb = -4.962997438e-02 lpdiblcb = 2.461187135e-8
+ drout = 1.009513028e+00 ldrout = -1.911563762e-8
+ pscbe1 = 8.087328239e+08 lpscbe1 = -8.726405225e+0
+ pscbe2 = 9.337822739e-09 lpscbe2 = -5.006721217e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.452507416e+00 lbeta0 = 4.140626236e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.281302899e+09 lbgidl = -4.276314530e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.536677683e-01 lkt1 = -1.884836796e-8
+ kt2 = -2.715603810e-02 lkt2 = -1.020745390e-8
+ at = 1.702205398e+05 lat = -6.751088280e-2
+ ute = 1.997060000e-02 lute = -1.995592161e-8
+ ua1 = 2.656528384e-09 lua1 = -2.522428491e-16
+ ub1 = -1.042863932e-18 lub1 = -3.149044430e-25
+ uc1 = -1.224595845e-10 luc1 = 2.607540497e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.42 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.415625649e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.875991477e-07 wvth0 = 7.712833416e-07 pvth0 = -3.850747776e-13
+ k1 = 1.983997073e+00 lk1 = -7.064144437e-07 wk1 = -3.081762099e-06 pk1 = 1.538615955e-12
+ k2 = -5.341717433e-01 lk2 = 2.574963977e-07 wk2 = 1.112814629e-06 pk2 = -5.555893956e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.286530863e+00 ldsub = -1.430548313e-07 wdsub = 2.557401725e-07 pdsub = -1.276821172e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-4.498653912e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.091290947e-07 wvoff = 4.481196497e-07 pvoff = -2.237304569e-13
+ nfactor = {1.884975111e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.218057618e-08 wnfactor = -7.105361633e-07 pnfactor = 3.547458376e-13
+ eta0 = -3.356492968e-01 leta0 = 2.058054720e-07 peta0 = -1.110223025e-28
+ etab = -3.749470590e-04 letab = -6.232944635e-11
+ u0 = -3.462248221e-03 lu0 = 5.614458706e-09 wu0 = 2.485866036e-08 pu0 = -1.241105907e-14
+ ua = -4.156515641e-09 lua = 1.481931175e-15 wua = 6.176354973e-15 pua = -3.083637866e-21
+ ub = 3.325258140e-18 lub = -9.695365530e-25 wub = -3.749934273e-24 pub = 1.872210935e-30
+ uc = 1.519759822e-11 luc = -2.354621073e-17 wuc = -1.206905973e-16 puc = 6.025659106e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.126339524e+05 lvsat = -1.106785392e-01 wvsat = -3.956271029e-01 pvsat = 1.975227655e-7
+ a0 = 1.489275913e+00 la0 = -1.541610062e-07 wa0 = 1.917591505e-07 pa0 = -9.573863226e-14
+ ags = -5.135474311e+00 lags = 3.189491700e-06 wags = 1.090549355e-05 pags = -5.444731238e-12
+ a1 = 0.0
+ a2 = 4.703575340e-01 la2 = 2.644269531e-07 wa2 = 1.477251346e-06 pa2 = -7.375398935e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.740979208e-02 lketa = 5.216216915e-09 wketa = 6.221399104e-08 pketa = -3.106126824e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.291500842e+00 lpclm = -2.904850491e-07 wpclm = -1.035333468e-06 ppclm = 5.169057641e-13
+ pdiblc1 = 2.068740150e+00 lpdiblc1 = -5.335845508e-07 wpdiblc1 = -9.075185981e-07 ppdiblc1 = 4.530922729e-13
+ pdiblc2 = 3.944086101e-03 lpdiblc2 = -1.461113202e-09 wpdiblc2 = -2.007020820e-08 ppdiblc2 = 1.002035250e-14
+ pdiblcb = -1.037009891e+00 lpdiblcb = 5.175761055e-07 wpdiblcb = 2.150463812e-06 ppdiblcb = -1.073651315e-12
+ drout = 2.810409167e+00 ldrout = -9.182400483e-07 wdrout = -2.650269320e-06 pdrout = 1.323186712e-12
+ pscbe1 = 7.834646021e+08 lpscbe1 = 3.889133508e+00 wpscbe1 = -1.587297278e+00 ppscbe1 = 7.924819757e-7
+ pscbe2 = 1.028651919e-08 lpscbe2 = -5.237181436e-16 wpscbe2 = -1.930140303e-15 ppscbe2 = 9.636514982e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.106539599e+01 lbeta0 = -8.904611877e-07 wbeta0 = -2.472571162e-06 pbeta0 = 1.234468241e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.272564884e-09 lagidl = -5.854206066e-16 wagidl = -2.375982295e-15 pagidl = 1.186244800e-21
+ bgidl = 1.139114877e+09 lbgidl = 2.822635763e+01 wbgidl = 4.293274392e+02 pbgidl = -2.143481639e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.371143572e-01 lkt1 = 7.274009322e-08 wkt1 = 2.902137045e-07 pkt1 = -1.448935452e-13
+ kt2 = -3.939003267e-02 lkt2 = -4.099448602e-09 wkt2 = -1.198423007e-08 pkt2 = 5.983306625e-15
+ at = -1.546231263e+05 lat = 9.467219016e-02 wat = 3.663090965e-01 pat = -1.828853110e-7
+ ute = -1.462721607e-01 lute = 6.304327033e-08 wute = 2.154597017e-07 pute = -1.075714880e-13
+ ua1 = -2.406752952e-09 lua1 = 2.275676307e-15 wua1 = 9.985605734e-15 pua1 = -4.985463447e-21
+ ub1 = 3.280044765e-18 lub1 = -2.473181454e-24 wub1 = -1.050158872e-23 pub1 = 5.243075691e-30
+ uc1 = 4.611635663e-10 luc1 = -2.653072074e-16 wuc1 = -9.815343010e-16 puc1 = 4.900457228e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.43 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {4.979821655e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.893963042e-07 wvth0 = -2.754583363e-06 pvth0 = 4.938003866e-13
+ k1 = -5.488912135e+00 lk1 = 1.156320270e-06 wk1 = 1.100629321e-05 pk1 = -1.973043153e-12
+ k2 = 2.173950218e+00 lk2 = -4.175436229e-07 wk2 = -3.974337960e-06 pk2 = 7.124596944e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.097585205e+00 ldsub = -9.595729190e-08 wdsub = -9.133577590e-07 pdsub = 1.637330787e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {6.624843524e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.681407642e-07 wvoff = -1.600427320e-06 pvoff = 2.869006036e-13
+ nfactor = {1.024755921e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.666031127e-07 wnfactor = 2.537629155e-06 pnfactor = -4.549080904e-13
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 5.648108911e-02 lu0 = -9.327317273e-09 wu0 = -8.878092986e-08 pu0 = 1.591531339e-14
+ ua = 1.108584089e-08 lua = -2.317454826e-15 wua = -2.205841062e-14 pua = 3.954300980e-21
+ ub = -6.209030164e-18 lub = 1.407027821e-24 wub = 1.339262240e-23 pub = -2.400828455e-30
+ uc = -2.609382890e-10 luc = 4.528480121e-17 wuc = 4.310378475e-16 puc = -7.726999973e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.269157846e+05 lvsat = 1.484448260e-01 wvsat = 1.412953939e+00 pvsat = -2.532931879e-7
+ a0 = 1.159465112e+00 la0 = -7.195071700e-08 wa0 = -6.848541089e-07 pa0 = 1.227703718e-13
+ ags = 2.407594930e+01 lags = -4.091893807e-06 wags = -3.894819125e-05 pags = 6.982047505e-12
+ a1 = 0.0
+ a2 = 3.754863313e+00 la2 = -5.542853798e-07 wa2 = -5.275897666e-06 pa2 = 9.457837950e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.716616948e-02 lketa = -2.334356015e-08 wketa = -2.221928251e-07 pketa = 3.983139680e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.432333858e+00 lpclm = 3.884716072e-07 wpclm = 3.697619530e-06 ppclm = -6.628537651e-13
+ pdiblc1 = -1.437962476e+00 lpdiblc1 = 3.405136791e-07 wpdiblc1 = 3.241137850e-06 ppdiblc1 = -5.810225767e-13
+ pdiblc2 = -3.212891336e-02 lpdiblc2 = 7.530623007e-09 wpdiblc2 = 7.167931501e-08 ppdiblc2 = -1.284959241e-14
+ pdiblcb = 4.276452586e+00 lpdiblcb = -8.068841188e-07 wpdiblcb = -7.680227900e-06 ppdiblcb = 1.376796055e-12
+ drout = -4.862782773e+00 ldrout = 9.944181405e-07 wdrout = 9.465247573e-06 pdrout = -1.696787606e-12
+ pscbe1 = 7.966776780e+08 lpscbe1 = 5.955761537e-01 wpscbe1 = 5.668918852e+00 ppscbe1 = -1.016238738e-6
+ pscbe2 = 5.280065017e-09 lpscbe2 = 7.242156546e-16 wpscbe2 = 6.893358224e-15 ppscbe2 = -1.235737862e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.771132884e+00 lbeta0 = 9.277433044e-07 wbeta0 = 8.830611291e-06 pbeta0 = -1.583019533e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.652544603e-09 lagidl = 8.915018097e-16 wagidl = 8.485651052e-15 pagidl = -1.521180236e-21
+ bgidl = 1.898611884e+09 lbgidl = -1.610896638e+02 wbgidl = -1.533312283e+03 pbgidl = 2.748692264e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 9.155728460e-02 lkt1 = -1.088922436e-07 wkt1 = -1.036477516e-06 pkt1 = 1.858041419e-13
+ kt2 = -7.387581867e-02 lkt2 = 4.496650845e-09 wkt2 = 4.280082167e-08 pkt2 = -7.672689297e-15
+ at = 7.765805717e+05 lat = -1.374442996e-01 wat = -1.308246773e+00 pat = 2.345228578e-7
+ ute = 4.309720005e-01 lute = -8.084349552e-08 wute = -7.694989346e-07 pute = 1.379442265e-13
+ ua1 = 2.175394081e-08 lua1 = -3.746739024e-15 wua1 = -3.566287762e-14 pua1 = 6.393105757e-21
+ ub1 = -2.244969874e-17 lub1 = 3.940343060e-24 wub1 = 3.750567399e-23 pub1 = -6.723454648e-30
+ uc1 = -2.080679910e-09 luc1 = 3.682854067e-16 wuc1 = 3.505479646e-15 puc1 = -6.284098088e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.44 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-1.269050275e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.996638185e-08 wvth0 = 3.598864257e-07 pvth0 = -7.063310933e-14
+ k1 = 3.690739784e-01 lk1 = 1.162584122e-07 wk1 = -1.939438274e-07 pk1 = 3.806438528e-14
+ k2 = 1.126493342e-01 lk2 = -5.257876565e-08 wk2 = 9.837868032e-08 pk2 = -1.930829169e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.181454340e+00 ldsub = -3.177826582e-07 wdsub = -2.432391268e-07 pdsub = 4.773932721e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.932586765e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.493071303e-09 wvoff = 6.366758970e-07 pvoff = -1.249571949e-13
+ nfactor = {1.609274304e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.665432960e-06 wnfactor = -3.008817794e-05 pnfactor = 5.905256243e-12
+ eta0 = -1.572766027e-02 leta0 = 9.925663924e-08 weta0 = 4.057114549e-06 peta0 = -7.962695869e-13
+ etab = -1.330653680e+00 letab = 2.610380788e-07 wetab = 2.693014686e-06 petab = -5.285445274e-13
+ u0 = 3.764136752e-02 lu0 = -6.514264426e-09 wu0 = -5.281569289e-08 pu0 = 1.036587196e-14
+ ua = 1.112548059e-08 lua = -2.545002831e-15 wua = -2.174341162e-14 pua = 4.267470681e-21
+ ub = -7.715009635e-18 lub = 1.836029685e-24 wub = 1.619997916e-23 pub = -3.179488909e-30
+ uc = -5.996019784e-11 luc = 1.013426964e-17 wuc = 1.212730211e-16 puc = -2.380164948e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.283925993e+05 lvsat = -1.231040027e-01 wvsat = -8.501769339e-01 pvsat = 1.668599759e-7
+ a0 = -7.327031787e+00 la0 = 1.586828390e-06 wa0 = 1.478539743e-05 pa0 = -2.901856026e-12
+ ags = 1.249999822e+00 lags = 2.967322565e-14
+ a1 = 0.0
+ a2 = -1.724821846e+00 la2 = 4.686212176e-07 wa2 = 3.735646070e-06 pa2 = -7.331765758e-13
+ b0 = 6.227509746e-23 lb0 = -1.222242200e-29 wb0 = -1.261887773e-28 pb0 = 2.476644037e-35
+ b1 = 0.0
+ keta = -6.291107170e-01 lketa = 1.091348641e-07 wketa = 4.258182338e-07 pketa = -8.357321565e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.444016295e+00 lpclm = -3.354808429e-07 wpclm = -2.272650383e-06 ppclm = 4.460417273e-13
+ pdiblc1 = 2.303137957e+00 lpdiblc1 = -3.614419153e-07 wpdiblc1 = -3.482697043e-07 ppdiblc1 = 6.835315351e-14
+ pdiblc2 = 6.018594809e-02 lpdiblc2 = -9.873411690e-09 wpdiblc2 = -3.032559695e-08 ppdiblc2 = 5.951853286e-15
+ pdiblcb = 3.628864403e+01 lpdiblcb = -7.166275044e-06 wpdiblcb = -6.371788587e-05 ppdiblcb = 1.250559087e-11
+ drout = -1.064617429e+00 ldrout = 3.432735561e-07 wdrout = -3.459889385e-12 pdrout = 6.790551907e-19
+ pscbe1 = 7.889611196e+08 lpscbe1 = 2.166545971e+00 wpscbe1 = 2.236822278e+01 ppscbe1 = -4.390099244e-6
+ pscbe2 = -3.593804523e-08 lpscbe2 = 8.882566645e-15 wpscbe2 = 9.193013794e-14 ppscbe2 = -1.804266852e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.034329304e+01 lbeta0 = -2.236812259e-06 wbeta0 = -1.290867800e-05 pbeta0 = 2.533521687e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.731440797e-08 lagidl = -3.335299528e-15 wagidl = -3.230632357e-14 pagidl = 6.340600596e-21
+ bgidl = 9.999998390e+08 lbgidl = 2.676576519e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.684936357e-01 lkt1 = 1.032621659e-08 wkt1 = 3.592903232e-07 pkt1 = -7.051611528e-14
+ kt2 = -2.468902279e-02 lkt2 = -4.730570723e-09 wkt2 = -1.553932845e-13 pkt2 = 3.049826292e-20
+ at = 1.897987439e+05 lat = -3.531363718e-02 wat = -4.904316368e-01 pat = 9.625456519e-8
+ ute = 1.415420638e+00 lute = -2.817228313e-07 wute = 9.114898096e-13 pute = -1.788935469e-19
+ ua1 = 5.039621037e-09 lua1 = -8.216125862e-16 wua1 = -3.592905901e-15 pua1 = 7.051616767e-22
+ ub1 = -2.283656623e-18 lub1 = 3.561241326e-25 wub1 = 1.590392439e-30 pub1 = -3.121383719e-37
+ uc1 = -8.009134101e-10 luc1 = 1.520371561e-16 wuc1 = 1.568901422e-15 puc1 = -3.079204376e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.45 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.103465450e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.372432872e-7
+ k1 = 4.212539000e-01 lk1 = 1.292480499e-6
+ k2 = 3.746785924e-02 lk2 = -5.455876137e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.342036093e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.900477982e-8
+ nfactor = {1.372957310e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.456178280e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.406882844e-02 lu0 = -3.649697542e-8
+ ua = -4.675899092e-10 lua = -2.058989945e-15
+ ub = 1.518950173e-18 lub = -2.543513577e-24 wub = -2.465190329e-38
+ uc = -7.214574862e-11 luc = -7.411055910e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.663233076e+00 la0 = -1.425397138e-6
+ ags = 5.586589101e-01 lags = -6.867219644e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.480543051e-02 lketa = 4.713717867e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.042871993e-01 lpclm = -2.882714742e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.362379205e-04 lpdiblc2 = 3.014921787e-9
+ pdiblcb = -3.449004373e-03 lpdiblcb = 3.837222522e-8
+ drout = 0.56
+ pscbe1 = 7.008645946e+08 lpscbe1 = 1.787834404e+3
+ pscbe2 = 9.666011755e-09 lpscbe2 = -6.109300570e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.681808713e-10 lalpha0 = -9.363273314e-15
+ alpha1 = -2.465499712e-11 lalpha1 = 2.493008321e-15 walpha1 = 1.809457590e-31 palpha1 = -4.549493369e-36
+ beta0 = 3.268475902e+00 lbeta0 = -5.369320704e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.851746450e-11 lagidl = 1.148245110e-15
+ bgidl = 1.563007487e+09 lbgidl = -1.125973593e+4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.257277191e-01 lkt1 = -5.962237055e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.559898067e-01 lute = 5.259768035e-7
+ ua1 = 2.139727641e-09 lua1 = 7.187183033e-15
+ ub1 = -7.305069847e-19 lub1 = -1.900516184e-23
+ uc1 = 4.334531165e-11 luc1 = 7.650412604e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.46 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.09160285+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4858803
+ k2 = 0.010187476
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.23615392+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4457689+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0122439126
+ ua = -5.7054319e-10
+ ub = 1.39176982e-18
+ uc = -1.0920239e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.5919606
+ ags = 0.52432155
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.031235975
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.060146165
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 790259600.0
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.4593183e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.45554
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.47 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.096965714e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.289897344e-8
+ k1 = 4.522097581e-01 lk1 = 2.693395874e-7
+ k2 = 2.269705454e-02 lk2 = -1.000674338e-07 pk2 = -8.881784197e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.356936746e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.681625035e-9
+ nfactor = {1.558435894e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.012531388e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.492833185e-02 lu0 = -2.147338093e-8
+ ua = -9.089350183e-11 lua = -3.836844963e-15
+ ub = 1.293690895e-18 lub = 7.845593095e-25
+ uc = -1.424170877e-10 luc = 2.656931686e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.214167700e+05 lvsat = -4.887892486e-01 wvsat = -3.725290298e-15
+ a0 = 1.651852193e+00 la0 = -4.790887229e-7
+ ags = 4.986878111e-01 lags = 2.050510707e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.745180763e-02 lketa = 4.972209241e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.124149426e-01 lpclm = 4.580068028e-06 ppclm = -1.421085472e-26
+ pdiblc1 = 0.39
+ pdiblc2 = 3.589658719e-04 lpdiblc2 = -5.757576728e-10
+ pdiblcb = -4.431168108e-04 lpdiblcb = -8.696847218e-9
+ drout = 0.56
+ pscbe1 = 7.805209898e+08 lpscbe1 = 7.790172373e+1
+ pscbe2 = 9.152466940e-09 lpscbe2 = 1.664395553e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -6.915519527e-01 lbeta0 = 2.952970233e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.918552200e-10 lagidl = -3.673533665e-16
+ bgidl = 8.017422366e+08 lbgidl = 1.585916388e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.102799397e-01 lkt1 = 4.378792836e-7
+ kt2 = -3.137221091e-02 lkt2 = -5.270546994e-8
+ at = -1.793770334e+05 lat = 1.434884425e+0
+ ute = 1.630094498e-01 lute = -3.941233465e-6
+ ua1 = 5.335468721e-09 lua1 = -2.268886504e-14
+ ub1 = -4.231141289e-18 lub1 = 2.040085581e-23
+ uc1 = 7.910528872e-10 luc1 = -2.921114695e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.48 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.095938434e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.879060751e-8
+ k1 = 5.981645711e-01 lk1 = -3.143723879e-7
+ k2 = -3.088465745e-02 lk2 = 1.142200316e-07 wk2 = -1.665334537e-22 pk2 = -1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.473007613e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.273819047e-8
+ nfactor = {1.242240996e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.632940483e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.086841217e-03 lu0 = 5.887553094e-9
+ ua = -1.527435151e-09 lua = 1.908265777e-15
+ ub = 1.866108470e-18 lub = -1.504690264e-24
+ uc = -6.690246480e-11 luc = -3.630981963e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.449391836e+05 lvsat = -1.829351138e-1
+ a0 = 1.910452889e+00 la0 = -1.513301435e-6
+ ags = 7.538877290e-01 lags = -8.155610292e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.126732654e-02 lketa = 6.498136366e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.351940539e-01 lpclm = -1.209303965e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = 1.975631812e-02 lpdiblcb = -8.947974034e-08 wpdiblcb = 5.551115123e-23 ppdiblcb = -3.330669074e-28
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.675630966e-08 lpscbe2 = -2.874538651e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.560060825e+00 lbeta0 = 4.527846154e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.142724829e+09 lbgidl = 2.222366395e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.431844278e-01 lkt1 = -2.303799486e-7
+ kt2 = -4.015072270e-02 lkt2 = -1.759787501e-8
+ at = 2.750948889e+05 lat = -3.826692271e-1
+ ute = -1.644657739e+00 lute = 3.288106654e-6
+ ua1 = -3.289890404e-09 lua1 = 1.180623182e-14 wua1 = 2.646977960e-29 pua1 = 1.058791184e-34
+ ub1 = 3.182174067e-18 lub1 = -9.246956829e-24 pub1 = -4.930380658e-44
+ uc1 = 9.232922993e-11 luc1 = -1.267336281e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.49 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.087705784e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.233135855e-8
+ k1 = 4.322060899e-01 lk1 = 1.742259510e-8
+ k2 = 3.068207834e-02 lk2 = -8.868188432e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.898963481e-01 ldsub = 3.400822775e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.235009021e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.844034868e-9
+ nfactor = {1.145902819e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.558995947e-7
+ eta0 = -5.889335829e-02 leta0 = 2.776846300e-7
+ etab = 6.922211054e-01 letab = -1.523881978e-06 wetab = 5.329070518e-21 petab = -1.243449788e-26
+ u0 = 1.261063863e-02 lu0 = -3.156716733e-9
+ ua = -2.729587568e-10 lua = -5.997649717e-16
+ ub = 1.001375792e-18 lub = 2.241395141e-25
+ uc = -1.218261949e-10 luc = 7.349727172e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.024470420e+04 lvsat = 2.637689452e-2
+ a0 = 1.186919436e+00 la0 = -6.676632695e-8
+ ags = 8.181288894e-02 lags = 5.280946760e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.564960160e-03 lketa = -1.239492287e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.804209211e-02 lpclm = 5.843405517e-7
+ pdiblc1 = 4.090022531e-01 lpdiblc1 = -3.799053949e-8
+ pdiblc2 = 1.580250000e-07 lpdiblc2 = 4.295260411e-10
+ pdiblcb = -0.025
+ drout = 1.299330017e-01 ldrout = 8.598178973e-7
+ pscbe1 = 800000000.0
+ pscbe2 = -4.525975301e-09 lpscbe2 = 1.380354094e-14 ppscbe2 = 5.293955920e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.783523713e+00 lbeta0 = 2.081819624e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.269248399e+09 lbgidl = -3.071750489e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443138732e-01 lkt1 = -2.819538791e-8
+ kt2 = -6.052627731e-02 lkt2 = 2.313825818e-8
+ at = 6.473381100e+04 lat = 3.789831325e-2
+ ute = 0.0
+ ua1 = 2.826536098e-09 lua1 = -4.221256071e-16
+ ub1 = -1.527945722e-18 lub1 = 1.698208119e-25
+ uc1 = 1.541511415e-10 luc1 = -2.503320121e-16 wuc1 = -8.271806126e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.50 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.090803540e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.542683752e-8
+ k1 = 3.303703168e-01 lk1 = 1.191835189e-7
+ k2 = 6.197639260e-02 lk2 = -4.013950137e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.608541037e-01 ldsub = 2.691766759e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.254154280e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.930916229e-9
+ nfactor = {1.415355000e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.866454611e-7
+ eta0 = 3.612140650e-01 leta0 = -1.421140143e-7
+ etab = -1.663840256e+00 letab = 8.304476780e-7
+ u0 = 1.111754745e-02 lu0 = -1.664722981e-09 wu0 = -2.220446049e-22
+ ua = -5.585029939e-10 lua = -3.144306096e-16
+ ub = 1.068261686e-18 lub = 1.573027816e-25
+ uc = -6.456159825e-11 luc = 1.627476450e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.236673570e+04 lvsat = 2.425642272e-2
+ a0 = 1.059796782e+00 la0 = 6.026289207e-8
+ ags = -3.136337212e-02 lags = 6.411877525e-7
+ a1 = 0.0
+ a2 = 6.003039853e-01 la2 = 1.995492381e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.697697029e-02 lketa = -3.192249000e-08 pketa = 2.220446049e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.360771286e-01 lpclm = 8.667157091e-8
+ pdiblc1 = -2.571078061e-01 lpdiblc1 = 6.276299288e-7
+ pdiblc2 = -1.566939902e-04 lpdiblc2 = 5.862627701e-10
+ pdiblcb = -4.962997438e-02 lpdiblcb = 2.461187135e-8
+ drout = 1.009513028e+00 ldrout = -1.911563762e-8
+ pscbe1 = 8.087328239e+08 lpscbe1 = -8.726405225e+0
+ pscbe2 = 9.337822739e-09 lpscbe2 = -5.006721217e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.452507416e+00 lbeta0 = 4.140626236e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.281302899e+09 lbgidl = -4.276314530e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.536677683e-01 lkt1 = -1.884836796e-8
+ kt2 = -2.715603810e-02 lkt2 = -1.020745390e-8
+ at = 1.702205398e+05 lat = -6.751088280e-2
+ ute = 1.997060000e-02 lute = -1.995592161e-8
+ ua1 = 2.656528384e-09 lua1 = -2.522428491e-16
+ ub1 = -1.042863932e-18 lub1 = -3.149044430e-25
+ uc1 = -1.224595845e-10 luc1 = 2.607540497e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.51 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.636078809e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.807750323e-8
+ k1 = 1.779017642e-01 lk1 = 1.953057308e-7
+ k2 = 1.180036084e-01 lk2 = -6.811192927e-08 wk2 = 4.440892099e-22
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.436409767e+00 ldsub = -2.178841223e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.872407073e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.199021815e-8
+ nfactor = {1.468558791e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.600826700e-7
+ eta0 = -3.356492968e-01 leta0 = 2.058054720e-07 weta0 = -1.776356839e-21 peta0 = -1.332267630e-27
+ etab = -3.749470590e-04 letab = -6.232944635e-11
+ u0 = 1.110640063e-02 lu0 = -1.659157764e-09 wu0 = 2.220446049e-22
+ ua = -5.368054278e-10 lua = -3.252634449e-16
+ ub = 1.127574320e-18 lub = 1.276900591e-25
+ uc = -5.553424759e-11 luc = 1.176772427e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.077301317e+04 lvsat = 5.081512593e-3
+ a0 = 1.601658145e+00 la0 = -2.102695211e-07 wa0 = -2.842170943e-20
+ ags = 1.255791501e+00 lags = -1.443625346e-9
+ a1 = 0.0
+ a2 = 1.336114410e+00 la2 = -1.678151535e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.094870464e-02 lketa = -1.298752791e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.847340437e-01 lpclm = 1.245237620e-8
+ pdiblc1 = 1.536880444e+00 lpdiblc1 = -2.680456149e-7
+ pdiblc2 = -7.818245877e-03 lpdiblc2 = 4.411407473e-09 wpdiblc2 = -2.775557562e-23 ppdiblc2 = -1.387778781e-29
+ pdiblcb = 2.232894046e-01 lpdiblcb = -1.116472224e-07 wpdiblcb = 1.679212325e-21 ppdiblcb = -7.771561172e-28
+ drout = 1.257194209e+00 ldrout = -1.427741826e-7
+ pscbe1 = 7.825343518e+08 lpscbe1 = 4.353574932e+0
+ pscbe2 = 9.155342529e-09 lpscbe2 = 4.103876969e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.616322685e+00 lbeta0 = -1.669896063e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.199016140e-10 lagidl = 1.097891793e-16
+ bgidl = 1.390726211e+09 lbgidl = -9.739437524e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.670319194e-01 lkt1 = -1.217611504e-8
+ kt2 = -4.641350204e-02 lkt2 = -5.928761668e-10
+ at = 6.005572284e+04 lat = -1.250944546e-2
+ ute = -2.000000083e-02 lute = 4.156137656e-16
+ ua1 = 3.445404059e-09 lua1 = -6.461008633e-16 pua1 = -1.323488980e-35
+ ub1 = -2.874508868e-18 lub1 = 5.995717658e-25
+ uc1 = -1.140737297e-10 luc1 = 2.188864117e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.52 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.11636700562893+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.961428255393082
+ k2 = -0.155247466831761
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.562303405039308
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.275460947389937+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.5119570622327+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 0.0044502003490566
+ ua = -1.84169558459119e-9
+ ub = 1.63984061966667e-18
+ uc = -8.324553995283e-12
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 101158.998341202
+ a0 = 0.758099999261006
+ ags = 1.24999997272013
+ a1 = 0.0
+ a2 = 0.662874470440252
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0730519999606918
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.734690420259434
+ pdiblc1 = 0.461536473183962
+ pdiblc2 = 0.00987941513820755
+ pdiblcb = -0.224616327814465
+ drout = 0.684413503600629
+ pscbe1 = 800000000.518868
+ pscbe2 = 9.31998164677673e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.94639467130503
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.20550031084906e-10
+ bgidl = 999999975.393082
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.515879992940252
+ kt2 = -0.0487919994941038
+ at = 9870.39612421382
+ ute = -0.0199999991650943
+ ua1 = 8.53380055896226e-10
+ ub1 = -4.69150049528303e-19
+ uc1 = -2.62609955581761e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.53 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-1.058121566e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.143154118e-08 wvth0 = -2.376128828e-11 pvth0 = 4.663509230e-18
+ k1 = 2.554142313e-01 lk1 = 1.385658424e-07 wk1 = -4.837013762e-12 pk1 = 9.493364956e-19
+ k2 = 1.703066823e-01 lk2 = -6.389488508e-08 wk2 = -2.744673651e-12 pk2 = 5.386833735e-19
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.038883481e+00 ldsub = -2.898009885e-07 wdsub = 3.124091148e-11 pdsub = -6.131497493e-18
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {7.986543680e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.973813279e-08 wvoff = 9.745034134e-12 pvoff = -1.912609129e-18
+ nfactor = {-1.540806813e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.954157020e-07 wnfactor = 1.597801754e-10 pnfactor = -3.135925613e-17
+ eta0 = 2.361973800e+00 leta0 = -3.674029378e-07 weta0 = 1.401514288e-11 peta0 = -2.750682015e-18
+ etab = 2.476144294e-01 letab = -4.872071160e-08 wetab = -3.127308435e-12 petab = 6.137811892e-19
+ u0 = 6.688219202e-03 lu0 = -4.392447701e-10 wu0 = 3.553431638e-14 pu0 = -6.974142541e-21
+ ua = -1.617436322e-09 lua = -4.401424424e-17 wua = -1.958104148e-20 pua = 3.843073106e-27
+ ub = 1.779154414e-18 lub = -2.734242193e-26 wub = -2.689203732e-29 pub = 5.277965690e-36
+ uc = 1.111295255e-11 luc = -3.814902221e-18 wuc = 5.169838462e-23 puc = -1.014658369e-29
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.301390432e+05 lvsat = -2.531426851e-02 wvsat = -9.121199250e-07 pvsat = 1.790172178e-13
+ a0 = 1.338085238e+00 la0 = -1.138308028e-07 wa0 = 4.264561994e-12 pa0 = -8.369842703e-19
+ ags = 1.249999822e+00 lags = 2.967321677e-14
+ a1 = 0.0
+ a2 = 4.644782956e-01 la2 = 3.893822526e-08 wa2 = 1.696616675e-11 pa2 = -3.329864711e-18
+ b0 = -1.167893467e-23 lb0 = 2.292166113e-30 wb0 = -1.248083260e-34 pb0 = 2.449550607e-41
+ b1 = 0.0
+ keta = -3.795544285e-01 lketa = 6.015569915e-08 wketa = -2.655921257e-12 pketa = 5.212643845e-19
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.112110262e+00 lpclm = -7.407430517e-08 wpclm = -3.134408757e-12 ppclm = 6.151747272e-19
+ pdiblc1 = 2.099040335e+00 lpdiblc1 = -3.213846954e-07 wpdiblc1 = -1.548177966e-11 ppdiblc1 = 3.038531482e-18
+ pdiblc2 = 4.241323970e-02 lpdiblc2 = -6.385251077e-09 wpdiblc2 = 1.886547194e-13 ppdiblc2 = -3.702631868e-20
+ pdiblcb = -1.053815362e+00 lpdiblcb = 1.627427485e-07 wpdiblcb = 6.989266979e-13 ppdiblcb = -1.371748510e-19
+ drout = -1.064637350e+00 ldrout = 3.432774658e-07 wdrout = 3.053089074e-11 pdrout = -5.992145276e-18
+ pscbe1 = 8.020694396e+08 lpscbe1 = -4.061584545e-01 wpscbe1 = 1.339054565e-03 ppscbe1 = -2.628095398e-10
+ pscbe2 = 1.793839480e-08 lpscbe2 = -1.691492858e-15 wpscbe2 = 1.217907357e-19 ppscbe2 = -2.390325897e-26
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.277805658e+01 lbeta0 = -7.520211236e-07 wbeta0 = -2.422723628e-11 pbeta0 = 4.754958354e-18
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.619007551e-09 lagidl = 3.806672688e-16 wagidl = -9.471010914e-21 pagidl = 1.858827951e-27
+ bgidl = 9.999998390e+08 lbgidl = 2.676576233e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.579276349e-01 lkt1 = -3.100051955e-08 wkt1 = -9.707316622e-13 pkt1 = 1.905206588e-19
+ kt2 = -2.468991748e-02 lkt2 = -4.730395127e-09 wkt2 = 1.371227476e-12 pkt2 = -2.691239605e-19
+ at = -9.762196435e+04 lat = 2.109698813e-02 wat = -2.233237002e-06 pat = 4.383062600e-13
+ ute = 1.415425886e+00 lute = -2.817238613e-07 wute = -8.043203907e-12 pute = 1.578599411e-18
+ ua1 = 2.933961916e-09 lua1 = -4.083453988e-16 wua1 = 5.524848526e-21 pua1 = -1.084334402e-27
+ ub1 = -2.283647466e-18 lub1 = 3.561223354e-25 wub1 = -1.403400289e-29 pub1 = 2.754383581e-36
+ uc1 = 1.185543005e-10 luc1 = -2.842217409e-17 wuc1 = 2.633733071e-21 puc1 = -5.169096216e-28
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.54 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.121329107e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.106456477e-06 wvth0 = 2.994506259e-08 pvth0 = 2.252460039e-12
+ k1 = 1.764697158e-01 lk1 = 8.718470018e-06 wk1 = 4.103346655e-07 pk1 = -1.244827534e-11
+ k2 = 1.373569331e-01 lk2 = -3.336250437e-06 wk2 = -1.674452532e-07 pk2 = 4.678021578e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.168575632e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.258989873e-06 wvoff = -2.907738531e-08 pvoff = 2.045075652e-12
+ nfactor = {1.574964309e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.795635710e-05 wnfactor = -3.386267566e-07 pnfactor = 6.606770600e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.739268410e-02 lu0 = 1.126401350e-07 wu0 = -5.571819136e-09 pu0 = -2.500003279e-13
+ ua = -2.166088169e-10 lua = 8.221814676e-18 wua = -4.207226168e-16 pua = -3.465291879e-21
+ ub = 1.501017826e-18 lub = 3.280737229e-23 wub = 3.006020794e-26 pub = -5.925911420e-29
+ uc = 8.093417837e-11 luc = -6.271262188e-15 wuc = -2.566097186e-16 puc = 9.270267866e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.603104387e+05 lvsat = 2.061306529e-04 wvsat = 3.455418267e-06 pvsat = -3.455392870e-10
+ a0 = 1.665873862e+00 la0 = 1.711640139e-05 wa0 = -4.426780589e-09 pa0 = -3.108183937e-11
+ ags = 3.940367627e-01 lags = 2.483558888e-05 wags = 2.759580812e-07 pags = -4.278335594e-11
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.083301313e-01 lketa = -3.952074146e-07 wketa = 8.972409825e-08 pketa = 1.452657114e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.463308160e-01 lpclm = -1.905378731e-05 wpclm = -9.086342191e-07 ppclm = 2.710776301e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -3.343372555e-04 lpdiblc2 = 1.029493865e-08 wpdiblc2 = 7.888308145e-10 ppdiblc2 = -1.220357962e-14
+ pdiblcb = -1.364159747e-01 lpdiblcb = 1.282871031e-05 wpdiblcb = 2.228941279e-07 ppdiblcb = -2.144059722e-11
+ drout = 0.56
+ pscbe1 = 4.140098219e+08 lpscbe1 = 6.885435555e+03 wpscbe1 = 4.808580977e+02 ppscbe1 = -8.545169982e-3
+ pscbe2 = 7.428964237e-09 lpscbe2 = 2.981964269e-13 wpscbe2 = 3.749989598e-15 ppscbe2 = -5.101113426e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.112351828e-09 lalpha0 = -4.024555748e-14 walpha0 = -2.588512304e-15 palpha0 = 5.176834353e-20
+ alpha1 = -4.357965834e-10 lalpha1 = 1.071553786e-14 walpha1 = 6.892015748e-16 palpha1 = -1.378352493e-20
+ beta0 = 6.857263639e+00 lbeta0 = -2.934057082e-04 wbeta0 = -6.015927950e-06 pbeta0 = 4.828388527e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.458222054e-10 lagidl = -1.973147656e-14 wagidl = -9.606062475e-17 pagidl = 3.500092800e-20
+ bgidl = 3.419938991e+09 lbgidl = -4.839700116e+04 wbgidl = -3.112796563e+03 pbgidl = 6.225364335e-2
+ cgidl = 300.0
+ egidl = 7.476257567e-01 legidl = -6.476209966e-05 wegidl = -1.085622827e-06 pegidl = 1.085614848e-10
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.152227325e-01 lkt1 = -3.780406353e-06 wkt1 = -1.852408352e-07 pkt1 = 5.337683582e-12
+ kt2 = -4.983212847e-02 lkt2 = 1.187104121e-06 wkt2 = 1.989971510e-08 pkt2 = -1.989956884e-12
+ at = 0.0
+ ute = -2.799511237e-01 lute = -1.401727293e-05 wute = -1.274645568e-07 pute = 2.437902405e-11
+ ua1 = 3.967416702e-10 lua1 = 8.666091397e-14 wua1 = 2.921788299e-15 pua1 = -1.332227689e-19
+ ub1 = 3.199380436e-18 lub1 = -1.612477725e-22 wub1 = -6.587717441e-24 pub1 = 2.384429952e-28
+ uc1 = -1.576718520e-09 luc1 = 6.872043373e-14 wuc1 = 2.715732442e-15 puc1 = -1.023724092e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.55 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.176653964e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.425722036e-7
+ k1 = 6.124092374e-01 wk1 = -2.121019761e-7
+ k2 = -2.946171933e-02 wk2 = 6.646442193e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.798093703e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff = 7.318015527e-8
+ nfactor = {-3.229232929e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.964879947e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.302489784e-02 wu0 = -1.807229492e-8
+ ua = -2.161977111e-10 wua = -5.939935784e-16
+ ub = 3.141446727e-18 wub = -2.933004394e-24
+ uc = -2.326404549e-10 wuc = 2.069207095e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.603207456e+05 wvsat = -1.382218103e-5
+ a0 = 2.521725384e+00 wa0 = -1.558575864e-6
+ ags = 1.635861844e+00 wags = -1.863288333e-6
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.280912283e-01 wketa = 1.623596233e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -2.063935624e-01 wpclm = 4.468037435e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.804285945e-04 wpdiblc2 = 1.786294085e-10
+ pdiblcb = 5.050431147e-01 wpdiblcb = -8.491751318e-7
+ drout = 0.56
+ pscbe1 = 7.582942521e+08 wpscbe1 = 5.358389633e+1
+ pscbe2 = 2.233933354e-08 wpscbe2 = -2.175651490e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -7.813560922e+00 wbeta0 = 1.812690194e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.407878807e-10 wagidl = 1.654050092e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -2.490598231e+00 wegidl = 4.342650902e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.042499969e-01 wkt1 = 8.165315224e-8
+ kt2 = 9.525258983e-03 wkt2 = -7.960178577e-8
+ at = 0.0
+ ute = -9.808405280e-01 wute = 1.091531444e-6
+ ua1 = 4.729946614e-09 wua1 = -3.739594949e-15
+ ub1 = -4.863304494e-18 wub1 = 5.334870473e-24
+ uc1 = 1.859429445e-09 wuc1 = -2.403076137e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.56 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.186346122e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.753013816e-08 wvth0 = 1.498294500e-07 pvth0 = -5.805263700e-14
+ k1 = 4.409497056e-01 lk1 = 1.371550232e-06 wk1 = 1.887536112e-08 pk1 = -1.847648930e-12
+ k2 = 3.133915398e-02 lk2 = -4.863622979e-07 wk2 = -1.448685500e-08 pk2 = 6.475507162e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.992694473e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.556663125e-07 wvoff = 1.065728307e-07 pvoff = -2.671168599e-13
+ nfactor = {-1.144808225e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.574475373e-06 wnfactor = 4.531480555e-06 pnfactor = -1.253165341e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.631717432e-02 lu0 = -1.063284421e-07 wu0 = -3.585437331e-08 pu0 = 1.422435573e-13
+ ua = 2.107057236e-09 lua = -1.858433198e-14 wua = -3.684451197e-15 pua = 2.472138946e-20
+ ub = 2.617825851e-18 lub = 4.188582145e-24 wub = -2.219663315e-24 pub = -5.706204327e-30
+ uc = -3.784830685e-10 luc = 1.166633714e-15 wuc = 3.957202364e-16 puc = -1.510257448e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.053701554e+04 lvsat = 7.182038493e-01 wvsat = 2.529215430e-01 pvsat = -2.023297014e-6
+ a0 = 2.581153989e+00 la0 = -4.753851653e-07 wa0 = -1.557799753e-06 pa0 = -6.208317961e-15
+ ags = 1.707516594e+00 lags = -5.731853377e-07 wags = -2.026374195e-06 pags = 1.304567030e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.581973174e-01 lketa = 2.408265851e-07 wketa = 2.024071470e-07 pketa = -3.203507544e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -2.994426075e+00 lpclm = 2.230221090e-05 wpclm = 4.160625046e-06 ppclm = -2.970784076e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 6.118628000e-03 lpdiblc2 = -4.750123066e-08 wpdiblc2 = -9.654990741e-09 ppdiblc2 = 7.866173348e-14
+ pdiblcb = 8.188054114e-01 lpdiblcb = -2.509867758e-06 wpdiblcb = -1.373316139e-06 ppdiblcb = 4.192742812e-12
+ drout = 0.56
+ pscbe1 = -6.842780468e+08 lpscbe1 = 1.153951810e+04 wpscbe1 = 2.455460203e+03 ppscbe1 = -1.921324507e-2
+ pscbe2 = 9.534387893e-08 lpscbe2 = -5.839827048e-13 wpscbe2 = -1.444836982e-13 ppscbe2 = 9.817272621e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -1.434065146e+01 lbeta0 = 5.221192687e-05 wbeta0 = 2.288014929e-05 pbeta0 = -3.802248518e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.452641166e-09 lagidl = 4.894376573e-15 wagidl = 2.756689026e-15 pagidl = -8.820301038e-21
+ bgidl = 1.478413642e+08 lbgidl = 6.816642750e+03 wbgidl = 1.096141879e+03 pbgidl = -8.768329368e-3
+ cgidl = 300.0
+ egidl = -5.080720440e+00 legidl = 2.071907393e-05 wegidl = 8.684503842e-06 pegidl = -3.473163226e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.531665487e-01 lkt1 = 2.791075961e-06 wkt1 = 5.747849373e-07 pkt1 = -3.944691829e-12
+ kt2 = 2.484443076e-02 lkt2 = -1.225421146e-07 wkt2 = -9.423663103e-08 pkt2 = 1.170680055e-13
+ at = -4.719889202e+05 lat = 3.775564450e+00 wat = 4.905088172e-01 pat = -3.923710014e-6
+ ute = 1.243299654e+00 lute = -1.779148672e-05 wute = -1.810903433e-06 pute = 2.321734573e-11
+ ua1 = 2.102712726e-08 lua1 = -1.303654667e-13 wua1 = -2.630411551e-14 pua1 = 1.804995796e-19
+ ub1 = -2.087332141e-17 lub1 = 1.280683680e-22 wub1 = 2.789748624e-23 pub1 = -1.804843426e-28
+ uc1 = 3.438494081e-09 luc1 = -1.263135647e-14 wuc1 = -4.437937442e-15 puc1 = 1.627739482e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.57 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.203919252e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.478097425e-07 wvth0 = 1.810095411e-07 pvth0 = -1.827500843e-13
+ k1 = 1.110703949e+00 lk1 = -1.306974471e-06 wk1 = -8.591759090e-07 pk1 = 1.663910783e-12
+ k2 = -2.065738911e-01 lk2 = 4.651150164e-07 wk2 = 2.945099707e-07 pk2 = -5.882094738e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.248243378e-01 ldsub = 3.938573505e-06 wdsub = 1.650872855e-06 pdsub = -6.602278030e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.441080725e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.493864316e-08 wvoff = -5.351942534e-09 pvoff = 1.804999683e-13
+ nfactor = {2.351269602e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.407266320e-06 wnfactor = -1.859077961e-06 pnfactor = 1.302588359e-11
+ eta0 = -1.821133918e-01 leta0 = 1.048260914e-06 weta0 = 4.393838240e-07 peta0 = -1.757212349e-12
+ etab = 1.591472712e-01 letab = -9.164206614e-07 wetab = -3.841223204e-07 petab = 1.536206952e-12
+ u0 = 6.388936871e-03 lu0 = 1.336251048e-08 wu0 = 2.846217431e-09 pu0 = -1.253036076e-14
+ ua = -4.140132074e-09 lua = 6.399833571e-15 wua = 4.379695203e-15 pua = -7.529268991e-21
+ ub = 5.208040525e-18 lub = -6.170372744e-24 wub = -5.602120806e-24 pub = 7.821139531e-30
+ uc = -3.831773218e-11 luc = -1.937776094e-16 wuc = -4.791693032e-17 puc = 2.639651456e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.467316719e+05 lvsat = -7.862982729e-01 wvsat = -5.058983696e-01 pvsat = 1.011424904e-6
+ a0 = 4.041568910e+00 la0 = -6.315971443e-06 wa0 = -3.572415360e-06 pa0 = 8.050773367e-12
+ ags = 2.725599454e+00 lags = -4.644768484e-06 wags = -3.305204025e-06 pags = 6.418946408e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.986990011e-01 lketa = 4.028035512e-07 wketa = 2.639046053e-07 pketa = -5.662953869e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.829780705e+00 lpclm = -1.298813043e-05 wpclm = -8.204854338e-06 ppclm = 1.974498815e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -1.102166880e-02 lpdiblc2 = 2.104735842e-08 wpdiblc2 = 1.883616275e-08 ppdiblc2 = -3.528193948e-14
+ pdiblcb = 4.073668452e-01 lpdiblcb = -8.644159009e-07 wpdiblcb = -6.497561780e-07 ppdiblcb = 1.299034785e-12
+ drout = 0.56
+ pscbe1 = 3.576165074e+09 lpscbe1 = -5.499122956e+03 wpscbe1 = -4.653718827e+03 ppscbe1 = 9.218245800e-3
+ pscbe2 = -8.072512267e-08 lpscbe2 = 1.201638909e-13 wpscbe2 = 1.634092948e-13 ppscbe2 = -2.496184086e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -1.385075071e+01 lbeta0 = 5.025268394e-05 wbeta0 = 3.253857630e-05 pbeta0 = -7.664909428e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.576261683e-10 lagidl = 9.150479168e-16 wagidl = 9.347554375e-16 pagidl = -1.533905803e-21
+ bgidl = 1.613464985e+09 lbgidl = 9.552255017e+02 wbgidl = -7.891073712e+02 pbgidl = -1.228718025e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.131372385e-01 lkt1 = -1.073428955e-06 wkt1 = -7.649374852e-07 pkt1 = 1.413213165e-12
+ kt2 = 2.610367839e-02 lkt2 = -1.275781796e-07 wkt2 = -1.110630476e-07 pkt2 = 1.843613043e-13
+ at = 8.454888671e+05 lat = -1.493378353e+00 wat = -9.561582704e-01 pat = 1.861895036e-6
+ ute = -6.632621542e+00 lute = 1.370640927e-05 wute = 8.361383580e-06 pute = -1.746432569e-11
+ ua1 = -2.509287044e-08 lua1 = 5.408062585e-14 wua1 = 3.654859707e-14 pua1 = -7.086507400e-20
+ ub1 = 2.302883931e-17 lub1 = -4.750800681e-23 wub1 = -3.326920310e-23 pub1 = 6.413745722e-29
+ uc1 = 3.378260804e-10 luc1 = -2.309634634e-16 wuc1 = -4.115293163e-16 puc1 = 1.747217237e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.58 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.112285685e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.539004192e-08 wvth0 = 4.120358219e-08 pvth0 = 9.675907626e-14
+ k1 = 6.836297566e-01 lk1 = -4.531399864e-07 wk1 = -4.214645097e-07 pk1 = 7.888097022e-13
+ k2 = -5.494558913e-02 lk2 = 1.619698592e-07 wk2 = 1.435386865e-07 pk2 = -2.863778694e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.512964069e+00 ldsub = -1.934844034e-06 wdsub = -3.558923898e-06 pdsub = 3.813486276e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.655175870e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.213535015e-08 wvoff = 7.043307297e-08 pvoff = 2.898563931e-14
+ nfactor = {-2.558744598e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.409153220e-06 wnfactor = 6.210144920e-06 pnfactor = -3.106631290e-12
+ eta0 = 4.686440022e-01 leta0 = -2.527755675e-07 weta0 = -8.843172078e-07 peta0 = 8.892167945e-13
+ etab = 2.566601823e-01 letab = -1.111374812e-06 wetab = 7.301360022e-07 petab = -6.914907135e-13
+ u0 = 1.357682281e-02 lu0 = -1.007978298e-09 wu0 = -1.619626135e-09 pu0 = -3.601956024e-15
+ ua = -2.466618091e-10 lua = -1.384245258e-15 wua = -4.408188909e-17 pua = 1.315033718e-21
+ ub = 1.224496530e-18 lub = 1.793787340e-24 wub = -3.740199707e-25 pub = -2.631219487e-30
+ uc = -2.763770956e-10 luc = 2.821661438e-16 wuc = 2.590755293e-16 puc = -3.497941342e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.323592483e+04 lvsat = 1.532914943e-01 wvsat = 1.064133402e-01 pvsat = -2.127484666e-7
+ a0 = 6.514605825e-01 la0 = 4.617534826e-07 wa0 = 8.975961021e-07 pa0 = -8.859640989e-13
+ ags = -1.812615073e-01 lags = 1.166816895e-06 wags = 4.409947674e-07 pags = -1.070697720e-12
+ a1 = 0.0
+ a2 = 1.459129381e+00 la2 = -1.317774301e-06 wa2 = -1.104906490e-06 pa2 = 2.209000875e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.470845467e-02 lketa = -4.384715584e-08 wketa = -4.571875257e-08 pketa = 5.272375556e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.351135812e+00 lpclm = 1.368424629e-06 wpclm = 2.328695590e-06 ppclm = -1.314369548e-12
+ pdiblc1 = -6.851537383e-01 lpdiblc1 = 2.149517239e-06 wpdiblc1 = 1.834146818e-06 ppdiblc1 = -3.666945539e-12
+ pdiblc2 = -1.417562207e-03 lpdiblc2 = 1.846204249e-09 wpdiblc2 = 2.376541438e-09 ppdiblc2 = -2.374794680e-15
+ pdiblcb = -0.025
+ drout = 1.616277352e-01 ldrout = 7.964517260e-07 wdrout = -5.313026201e-08 pdrout = 1.062214733e-13
+ pscbe1 = 8.060215384e+08 lpscbe1 = 3.912805907e+01 wpscbe1 = -1.009397713e+01 ppscbe1 = -6.559083496e-5
+ pscbe2 = -5.087362719e-08 lpscbe2 = 6.048284079e-14 wpscbe2 = 7.769312504e-14 ppscbe2 = -7.824907049e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.750496186e+00 lbeta0 = 3.067537073e-06 wbeta0 = -4.973571560e-06 pbeta0 = -1.652369988e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.245084270e-09 lagidl = -2.489121468e-15 wagidl = -1.919518503e-15 pagidl = 4.172544186e-21
+ bgidl = 2.157293133e+09 lbgidl = -1.320310822e+02 wbgidl = -1.488640045e+03 pbgidl = 1.698331654e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.965922154e-01 lkt1 = -5.434469784e-08 wkt1 = -7.999638772e-08 pkt1 = 4.383440202e-14
+ kt2 = -7.492061447e-02 lkt2 = 7.439615328e-08 wkt2 = 2.412940011e-08 pkt2 = -8.592422465e-14
+ at = -4.039955183e+04 lat = 2.777473567e-01 wat = 1.762363177e-01 pat = -4.020618298e-7
+ ute = -3.008496165e+00 lute = 6.460822246e-06 wute = 5.043178223e-06 pute = -1.083035386e-11
+ ua1 = -7.830996148e-09 lua1 = 1.956956475e-14 wua1 = 1.786534919e-14 pua1 = -3.351231045e-20
+ ub1 = 7.314834016e-18 lub1 = -1.609154602e-23 wub1 = -1.482325779e-23 pub1 = 2.725912436e-29
+ uc1 = 1.078887165e-09 luc1 = -1.712540953e-15 wuc1 = -1.550146093e-15 puc1 = 2.451118394e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.59 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.179971196e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.224572083e-08 wvth0 = 1.494728123e-07 pvth0 = -1.143057593e-14
+ k1 = -2.830053748e-01 lk1 = 5.127846681e-07 wk1 = 1.028209032e-06 pk1 = -6.597983296e-13
+ k2 = 2.834346381e-01 lk2 = -1.761616585e-07 wk2 = -3.712331144e-07 pk2 = 2.280155742e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.274697401e+00 ldsub = 2.849298505e-06 wdsub = 4.585637814e-06 pdsub = -4.325089183e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.376290035e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.992306451e-08 wvoff = 1.881049633e-07 pvoff = -8.859976215e-14
+ nfactor = {1.151056629e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.627317611e-07 wnfactor = 2.179623566e-06 pnfactor = 9.209276300e-13
+ eta0 = 1.716185986e+00 leta0 = -1.499400608e-06 weta0 = -2.271355690e-06 peta0 = 2.275235804e-12
+ etab = -1.709719861e+00 letab = 8.535599425e-07 wetab = 7.690853273e-08 petab = -3.874336629e-14
+ u0 = 2.007586128e-02 lu0 = -7.502239981e-09 wu0 = -1.501692897e-08 pu0 = 9.785499797e-15
+ ua = -4.726996842e-10 lua = -1.158373521e-15 wua = -1.438331177e-16 pua = 1.414711629e-21
+ ub = 3.094534331e-18 lub = -7.487598286e-26 wub = -3.396665150e-24 pub = 3.892040490e-31
+ uc = 5.126249913e-11 luc = -4.523263585e-17 wuc = -1.941573243e-16 puc = 1.031055933e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.806678373e+04 lvsat = 8.204119326e-02 wvsat = -9.555058908e-03 pvsat = -9.686530429e-8
+ a0 = -4.814589115e-01 la0 = 1.593840281e-06 wa0 = 2.583625414e-06 pa0 = -2.570754179e-12
+ ags = 7.107681688e-01 lags = 2.754428605e-07 wags = -1.244044008e-06 pags = 6.131025513e-13
+ a1 = 0.0
+ a2 = -7.505600368e-01 la2 = 8.902909945e-07 wa2 = 2.264469571e-06 pa2 = -1.157898695e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.902331606e-02 lketa = -5.815149580e-08 wketa = -3.695655397e-08 pketa = 4.396799717e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -2.917597307e+00 lpclm = 2.933734775e-06 wpclm = 5.789435900e-06 ppclm = -4.772566214e-12
+ pdiblc1 = -1.325955106e+00 lpdiblc1 = 2.789847618e-06 wpdiblc1 = 1.791721556e-06 ppdiblc1 = -3.624551459e-12
+ pdiblc2 = -3.375724211e-03 lpdiblc2 = 3.802927004e-09 wpdiblc2 = 5.396098988e-09 ppdiblc2 = -5.392132855e-15
+ pdiblcb = -1.128478045e-01 lpdiblcb = 8.778323634e-08 wpdiblcb = 1.059728072e-07 ppdiblcb = -1.058949172e-13
+ drout = 1.040889238e+00 ldrout = -8.216351981e-08 wdrout = -5.259631778e-08 pdrout = 1.056879215e-13
+ pscbe1 = 9.278260803e+08 lpscbe1 = -8.258695646e+01 wpscbe1 = -1.996374549e+02 ppscbe1 = 1.238133284e-4
+ pscbe2 = 1.036766058e-08 lpscbe2 = -7.134346404e-16 wpscbe2 = -1.726329532e-15 ppscbe2 = 1.112010780e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.460711488e+01 lbeta0 = -1.785512005e-06 wbeta0 = -1.031704234e-05 pbeta0 = 3.687173345e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.284889185e-09 lagidl = 1.038257456e-15 wagidl = 3.997818359e-15 pagidl = -1.740443433e-21
+ bgidl = 2.209106220e+09 lbgidl = -1.838060862e+02 wbgidl = -1.555287840e+03 pbgidl = 2.364319744e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.642297497e-01 lkt1 = 1.131696229e-07 wkt1 = 1.853363762e-07 pkt1 = -2.213033423e-13
+ kt2 = 9.578227301e-02 lkt2 = -9.618126758e-08 wkt2 = -2.060829662e-07 pkt2 = 1.441189356e-13
+ at = 4.401061454e+05 lat = -2.024051688e-01 wat = -4.524124794e-01 pat = 2.261249104e-7
+ ute = 6.341010916e+00 lute = -2.881812947e-06 wute = -1.059603573e-05 pute = 4.797365273e-12
+ ua1 = 2.270792566e-08 lua1 = -1.094691096e-14 wua1 = -3.361239788e-14 pua1 = 1.792760048e-20
+ ub1 = -1.841247844e-17 lub1 = 9.616856862e-24 wub1 = 2.911689324e-23 pub1 = -1.664873066e-29
+ uc1 = -1.610760969e-09 luc1 = 9.751302899e-16 wuc1 = 2.494857471e-15 puc1 = -1.590912092e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.60 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-7.863276756e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.642867115e-07 wvth0 = -2.971769354e-07 pvth0 = 2.115660104e-13
+ k1 = -8.705093437e-01 lk1 = 8.061048372e-07 wk1 = 1.757464121e-06 pk1 = -1.023889872e-12
+ k2 = 5.487550268e-01 lk2 = -3.086268424e-07 wk2 = -7.220737716e-07 pk2 = 4.031780350e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.121749607e+00 ldsub = -1.842018611e-06 wdsub = -9.530403398e-06 pdsub = 2.722556133e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-5.266849074e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.234774591e-08 wvoff = -2.255850215e-07 pvoff = 1.179411681e-13
+ nfactor = {-2.995410550e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.290240116e-06 wnfactor = 7.483005374e-06 pnfactor = -1.726865288e-12
+ eta0 = -3.058835446e+00 leta0 = 8.846004675e-07 weta0 = 4.564909620e-06 peta0 = -1.137872196e-12
+ etab = 2.484570086e-03 letab = -1.283802877e-09 wetab = -4.793442904e-09 petab = 2.047570569e-15
+ u0 = 1.472627811e-02 lu0 = -4.831380339e-09 wu0 = -6.068044059e-09 pu0 = 5.317634771e-15
+ ua = -1.695792232e-09 lua = -5.477262195e-16 wua = 1.942823488e-15 pua = 3.729170185e-22
+ ub = 3.927024256e-18 lub = -4.905090650e-25 wub = -4.692751520e-24 pub = 1.036294610e-30
+ uc = -4.272392067e-11 luc = 1.691494027e-18 wuc = -2.147410474e-17 puc = 1.689090568e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.796598136e+05 lvsat = -3.358510081e-02 wvsat = -3.333963302e-01 pvsat = 6.481730805e-8
+ a0 = 4.115378657e+00 la0 = -7.011998281e-07 wa0 = -4.213779860e-06 pa0 = 8.229523648e-13
+ ags = 2.187791688e+00 lags = -4.619832868e-07 wags = -1.562323097e-06 pags = 7.720081609e-13
+ a1 = 0.0
+ a2 = 1.852267595e+00 la2 = -4.092097429e-07 wa2 = -8.652337775e-07 pa2 = 4.046526470e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.884969050e-02 lketa = -6.305746064e-08 wketa = -1.170038873e-07 pketa = 8.393282907e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.859735891e+00 lpclm = -9.492154839e-07 wpclm = -6.998605697e-06 ppclm = 1.612055374e-12
+ pdiblc1 = 7.877757338e+00 lpdiblc1 = -1.805243876e-06 wpdiblc1 = -1.062928803e-05 ppdiblc1 = 2.576823891e-12
+ pdiblc2 = -3.636146721e-03 lpdiblc2 = 3.932946848e-09 wpdiblc2 = -7.010503001e-09 ppdiblc2 = 8.020492868e-16
+ pdiblcb = 3.764576247e-01 lpdiblcb = -1.565098387e-07 wpdiblcb = -2.567577254e-07 ppdiblcb = 7.520374216e-14
+ drout = 4.252533759e-01 ldrout = 2.252019190e-07 wdrout = 1.394592402e-06 pdrout = -6.168427548e-13
+ pscbe1 = 7.248333207e+08 lpscbe1 = 1.876022369e+01 wpscbe1 = 9.672493090e+01 ppscbe1 = -2.415003818e-5
+ pscbe2 = 8.015599920e-09 lpscbe2 = 4.608669252e-16 wpscbe2 = 1.910564213e-15 ppscbe2 = -7.037629750e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.314296727e+01 lbeta0 = -1.054514348e-06 wbeta0 = -5.911756633e-06 pbeta0 = 1.487768375e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.454925981e-09 lagidl = 6.238858774e-16 wagidl = 2.237917366e-15 pagidl = -8.617864642e-22
+ bgidl = 3.535663444e+09 lbgidl = -8.461096785e+02 wbgidl = -3.595584021e+03 pbgidl = 1.255080447e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.647761481e-01 lkt1 = -8.626357951e-08 wkt1 = -5.066749766e-07 pkt1 = 1.241937057e-13
+ kt2 = -1.585777298e-01 lkt2 = 3.081177920e-08 wkt2 = 1.880222409e-07 pkt2 = -5.264400065e-14
+ at = 2.639605941e+05 lat = -1.144618601e-01 wat = -3.418081826e-01 pat = 1.709040562e-7
+ ute = -1.619851232e+00 lute = 1.092766894e-06 wute = 2.681849817e-06 pute = -1.831818256e-12
+ ua1 = -1.140747603e-09 lua1 = 9.598969037e-16 wua1 = 7.687821066e-15 pua1 = -2.692153329e-21
+ ub1 = 3.135044707e-18 lub1 = -1.141067284e-24 wub1 = -1.007388677e-23 pub1 = 2.917854127e-30
+ uc1 = 4.554193161e-10 luc1 = -5.644121018e-17 wuc1 = -9.546480266e-16 puc1 = 1.313052698e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.61 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-2.236007191e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.105077672e-07 wvth0 = 1.876866278e-06 pvth0 = -3.528766963e-13
+ k1 = 7.384333277e+00 lk1 = -1.336894073e-06 wk1 = -1.076679276e-05 pk1 = 2.241051577e-12
+ k2 = -2.629105617e+00 lk2 = 5.164777140e-07 wk2 = 4.146958103e-06 pk2 = -8.657777897e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.483808842e+00 ldsub = 1.122508802e-06 wdsub = 8.458858513e-06 pdsub = -1.881674974e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.406094005e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.617239354e-07 wvoff = 1.895293762e-06 pvoff = -4.387309736e-13
+ nfactor = {4.099333271e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.108468144e-07 wnfactor = -2.660937788e-06 pnfactor = 8.563386452e-13
+ eta0 = -2.533352966e+00 leta0 = 8.050130775e-07 weta0 = 5.068082857e-06 peta0 = -1.349453082e-12
+ etab = -2.491714952e-01 letab = 6.563584335e-08 wetab = 4.166414725e-07 petab = -1.100261518e-13
+ u0 = -3.931520053e-02 lu0 = 9.228471372e-09 wu0 = 7.336446668e-08 pu0 = -1.546979730e-14
+ ua = -1.246469730e-08 lua = 2.282301080e-15 wua = 1.780746524e-14 pua = -3.825848688e-21
+ ub = 4.962086306e-18 lub = -7.995628301e-25 wub = -5.569120311e-24 pub = 1.340316767e-30
+ uc = -1.881996515e-10 luc = 4.054195026e-17 wuc = 3.015267845e-16 puc = -6.796095772e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -8.067986409e+04 lvsat = 6.007022249e-02 wvsat = 3.048186672e-01 pvsat = -1.006964348e-7
+ a0 = 1.910612541e+00 la0 = -1.619699637e-07 wa0 = -1.931970604e-06 pa0 = 2.715121939e-13
+ ags = -2.232709364e+00 lags = 6.835339303e-07 wags = 5.838107454e-06 pags = -1.145816130e-12
+ a1 = 0.0
+ a2 = -1.166886813e+00 la2 = 3.667770925e-07 wa2 = 3.067250797e-06 pa2 = -6.148328414e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.355870182e-01 lketa = 3.500402865e-08 wketa = 4.400906014e-07 pketa = -5.867767327e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.823378825e+00 lpclm = -2.054768492e-07 wpclm = -1.824981436e-06 ppclm = 3.444433080e-13
+ pdiblc1 = 4.100420548e-01 lpdiblc1 = 6.002878202e-08 wpdiblc1 = 8.632071141e-08 ppdiblc1 = -1.006269676e-13
+ pdiblc2 = -2.122074516e-04 lpdiblc2 = 3.289500638e-09 wpdiblc2 = 1.691670805e-08 ppdiblc2 = -5.514229393e-15
+ pdiblcb = -3.301491190e-01 lpdiblcb = 2.096075511e-08 wpdiblcb = 1.769058842e-07 ppdiblcb = -3.513676532e-14
+ drout = 2.644577102e+00 ldrout = -3.503674274e-07 wdrout = -3.285845763e-06 pdrout = 5.873251230e-13
+ pscbe1 = 8.003632026e+08 lpscbe1 = -7.128352767e-02 wpscbe1 = -6.088400677e-01 ppscbe1 = 1.194934328e-7
+ pscbe2 = 1.057066178e-08 lpscbe2 = -1.880252627e-16 wpscbe2 = -2.096530121e-15 ppscbe2 = 3.151890042e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.082389807e+00 lbeta0 = 1.286081894e-06 wbeta0 = 8.153589722e-06 pbeta0 = -2.155874512e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.536155632e-08 lagidl = -3.811205448e-15 wagidl = -2.521341933e-14 pagidl = 6.388769426e-21
+ bgidl = -2.266519172e+09 lbgidl = 6.411033646e+02 wbgidl = 5.475705246e+03 pbgidl = -1.074689263e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.602942008e-01 lkt1 = 6.641881472e-08 wkt1 = 4.097144696e-07 pkt1 = -1.113386561e-13
+ kt2 = -3.642300228e-02 lkt2 = 3.876297281e-10 wkt2 = -2.073429846e-08 pkt2 = -6.497883647e-16
+ at = -5.909520052e+05 lat = 1.053650859e-01 wat = 1.007165801e+00 pat = -1.766247579e-7
+ ute = 8.175024886e+00 lute = -1.440738537e-06 wute = -1.373741855e-05 pute = 2.415127298e-12
+ ua1 = 4.006223756e-09 lua1 = -3.450959675e-16 wua1 = -5.285149729e-15 pua1 = 5.784885114e-22
+ ub1 = -1.144613343e-18 lub1 = -7.936550384e-26 wub1 = 1.132287224e-24 pub1 = 1.330413465e-31
+ uc1 = 7.030159785e-10 luc1 = -1.262168548e-16 wuc1 = -1.222495743e-15 puc1 = 2.115788283e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.62 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-9.131464151e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.912350296e-08 wvth0 = -2.430473466e-07 pvth0 = 6.318815134e-14
+ k1 = -2.461972407e+00 lk1 = 5.955911123e-07 wk1 = 4.555182993e-06 pk1 = -7.661159949e-13
+ k2 = 1.401728314e+00 lk2 = -2.746339075e-07 wk2 = -2.064249603e-06 pk2 = 3.532648908e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.582313673e+00 ldsub = -1.245648734e-06 wdsub = -9.292487312e-06 pdsub = 1.602292914e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.454730825e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.997558499e-07 wvoff = -2.304693604e-06 pvoff = 3.855795468e-13
+ nfactor = {-1.592283436e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.418803916e-06 wnfactor = 2.410892514e-05 pnfactor = -4.397648502e-12
+ eta0 = 9.614531917e+00 leta0 = -1.579191549e-06 weta0 = -1.215753619e-05 peta0 = 2.031333040e-12
+ etab = 1.152236708e+00 letab = -2.094115378e-07 wetab = -1.516432309e-06 petab = 2.693685740e-13
+ u0 = 1.732488758e-02 lu0 = -1.887995521e-09 wu0 = -1.783033930e-08 pu0 = 2.428551295e-15
+ ua = 1.278425381e-10 lua = -1.891737506e-16 wua = -2.925651477e-15 pua = 2.433364654e-22
+ ub = 1.486926783e-18 lub = -1.175106462e-25 wub = 4.898377936e-25 pub = 1.511553543e-31
+ uc = 1.019148668e-10 luc = -1.639737569e-17 wuc = -1.522122869e-16 puc = 2.109214112e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.797713682e+05 lvsat = -1.088062386e-01 wvsat = -9.213561740e-01 pvsat = 1.399587704e-7
+ a0 = 3.578275269e+00 la0 = -4.892737889e-07 wa0 = -3.755253167e-06 pa0 = 6.293587460e-13
+ ags = 1.249999233e+00 lags = 1.275425170e-13 wags = 9.867348467e-13 pags = -1.640594691e-19
+ a1 = 0.0
+ a2 = -1.508118483e-01 la2 = 1.673571395e-07 wa2 = 1.031435218e-06 pa2 = -2.152734968e-13
+ b0 = -5.019913627e-23 lb0 = 9.852333480e-30 wb0 = 6.457175137e-29 pb0 = -1.267317478e-35
+ b1 = 0.0
+ keta = -1.474662724e+00 lketa = 2.585647221e-07 wketa = 1.835740521e-06 pketa = -3.325949048e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.398674527e+00 lpclm = -3.183872602e-07 wpclm = -2.156686251e-06 ppclm = 4.095453534e-13
+ pdiblc1 = 7.754236004e+00 lpdiblc1 = -1.381379443e-06 wpdiblc1 = -9.479887845e-06 ppdiblc1 = 1.776884955e-12
+ pdiblc2 = 1.563868345e-01 lpdiblc2 = -2.744541033e-08 wpdiblc2 = -1.910551160e-07 ppdiblc2 = 3.530336066e-14
+ pdiblcb = -3.787442150e+00 lpdiblcb = 6.995063719e-07 wpdiblcb = 4.582412087e-06 ppdiblcb = -8.997834402e-13
+ drout = -6.658353065e+00 ldrout = 1.475472162e-06 wdrout = 9.376843308e-06 pdrout = -1.897917547e-12
+ pscbe1 = 8.088983729e+08 lpscbe1 = -1.746438720e+00 wpscbe1 = -1.144608385e+01 ppscbe1 = 2.246465083e-6
+ pscbe2 = 4.665692959e-08 lpscbe2 = -7.270496615e-15 wpscbe2 = -4.814110270e-14 ppscbe2 = 9.352127041e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.710449712e+01 lbeta0 = -3.232351997e-06 wbeta0 = -2.401560842e-05 pbeta0 = 4.157813162e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.239381491e-08 lagidl = 1.636202486e-15 wagidl = 1.806192940e-14 pagidl = -2.104666892e-21
+ bgidl = 9.999993081e+08 lbgidl = 1.150455723e-04 wbgidl = 8.900520248e-04 pbgidl = -1.479844999e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.570337597e-01 lkt1 = -1.332470575e-07 wkt1 = -1.030868136e-06 pkt1 = 1.713972890e-13
+ kt2 = 6.915198019e-02 lkt2 = -2.033304421e-08 wkt2 = -1.573069279e-07 pkt2 = 2.615463876e-14
+ at = -5.161341296e+05 lat = 9.068095556e-02 wat = 7.015547315e-01 pat = -1.166440013e-7
+ ute = 7.004021545e+00 lute = -1.210911566e-06 wute = -9.368238009e-06 pute = 1.557610079e-12
+ ua1 = 1.119075317e-08 lua1 = -1.755167632e-15 wua1 = -1.384095273e-14 pua1 = 2.257693187e-21
+ ub1 = -9.348166561e-18 lub1 = 1.530704869e-24 wub1 = 1.184232410e-23 pub1 = -1.968964041e-30
+ uc1 = 6.823789804e-10 luc1 = -1.221665344e-16 wuc1 = -9.451434431e-16 puc1 = 1.571442791e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.63 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.000673396e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.302804208e-06 wvth0 = -1.252558272e-07 pvth0 = 2.505024481e-12
+ k1 = 1.050452350e+00 lk1 = -1.205825004e-05 wk1 = -7.138796846e-07 pk1 = 1.427706899e-11
+ k2 = -1.092550679e-01 lk2 = 2.629180932e-06 wk2 = 1.497747230e-07 pk2 = -2.995384376e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.090257148e-04 lcit = -1.980441513e-09 wcit = -1.273779653e-10 pcit = 2.547465683e-15
+ voff = {-2.192303752e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.019749918e-06 wvoff = -2.798240049e-07 pvoff = 5.596274427e-12
+ nfactor = {-4.187704613e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.233900155e-04 wnfactor = 7.073963429e-06 pnfactor = -1.414740692e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.082173069e-02 lu0 = -4.369145565e-07 wu0 = -2.284576291e-08 pu0 = 4.568984665e-13
+ ua = 1.979574033e-09 lua = -5.314908815e-14 wua = -3.245698970e-15 pua = 6.491159382e-20
+ ub = 3.081884836e-18 lub = -4.441044237e-23 wub = -2.003427997e-24 pub = 4.006708742e-29
+ uc = -1.547836563e-10 luc = 1.660073937e-15 wuc = 4.659696082e-17 puc = -9.319049677e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.807031471e+05 lvsat = -1.640725995e+01 wvsat = -1.055277530e+00 pvsat = 2.110477497e-5
+ a0 = 2.972090385e+00 la0 = -3.323932611e-05 wa0 = -1.684628769e-06 pa0 = 3.369133718e-11
+ ags = 4.815418726e+00 lags = -9.255875285e-05 wags = -5.411318594e-06 pags = 1.082223946e-10
+ a1 = 0.0
+ a2 = -9.399250686e-01 la2 = 3.479722253e-05 wa2 = 2.238086495e-06 pa2 = -4.476008490e-11
+ b0 = 1.327358130e-06 lb0 = -2.654618700e-11 wb0 = -1.707396691e-12 pb0 = 3.414667889e-17
+ b1 = -6.113584948e-09 lb1 = 1.222672055e-13 wb1 = 7.863977682e-15 pb1 = -1.572737736e-19
+ keta = -5.973718320e-01 lketa = 1.190959495e-05 wketa = 7.187843063e-07 pketa = -1.437515782e-11
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.020080816e-01 lpclm = -7.220716660e-06 wpclm = -5.943589540e-07 ppclm = 1.188674223e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -9.855324331e-03 lpdiblc2 = 2.034849687e-07 wpdiblc2 = 1.303579074e-08 ppdiblc2 = -2.607062335e-13
+ pdiblcb = 2.324044943e+00 lpdiblcb = -4.958146728e-05 wpdiblcb = -2.942026276e-06 ppdiblcb = 5.883836314e-11
+ drout = 0.56
+ pscbe1 = 6.881452110e+08 lpscbe1 = 2.236038602e+03 wpscbe1 = 1.282344570e+02 ppscbe1 = -2.564594888e-3
+ pscbe2 = 3.178954161e-09 lpscbe2 = 4.492852160e-14 wpscbe2 = 9.216828560e-15 ppscbe2 = -1.843297968e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.123485334e-09 lalpha0 = -2.046895443e-14 walpha0 = -1.316521468e-15 palpha0 = 2.632946171e-20
+ alpha1 = 1.123485334e-09 lalpha1 = -2.046895443e-14 walpha1 = -1.316521468e-15 palpha1 = 2.632946171e-20
+ beta0 = -2.741606575e+02 lbeta0 = 5.608578813e-03 wbeta0 = 3.554607962e-04 pbeta0 = -7.108954661e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.788412182e-08 lagidl = 3.665709191e-13 wagidl = 2.309607274e-14 pagidl = -4.619044792e-19
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -9.635519618e-02 legidl = 1.963537530e-05 pegidl = 7.105427358e-27
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.361926036e-01 lkt1 = 3.908278438e-06 wkt1 = 2.276265617e-07 pkt1 = -4.552363929e-12
+ kt2 = 1.763226918e-01 lkt2 = -4.573455196e-06 wkt2 = -2.710059441e-07 pkt2 = 5.419919693e-12
+ at = -7.265722389e+05 lat = 1.453091075e+01 wat = 9.345985898e-01 pat = -1.869128487e-5
+ ute = -2.904084825e+00 lute = 5.543433681e-05 wute = 3.247990113e-06 pute = -6.495741498e-11
+ ua1 = 6.853219243e-09 lua1 = -1.006062015e-13 wua1 = -5.383256281e-15 pua1 = 1.076611689e-19
+ ub1 = -6.547149141e-18 lub1 = 1.166209193e-22 wub1 = 5.949360512e-24 pub1 = -1.189828375e-28
+ uc1 = 5.198241713e-09 luc1 = -1.041362326e-13 wuc1 = -5.998980206e-15 puc1 = 1.199751949e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.64 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.065816+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44751769
+ k2 = 0.02220881
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.22291792+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9820229+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0089752
+ ua = -6.7797804e-10
+ ub = 8.6128111e-19
+ uc = -7.1776909e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160310.0
+ a0 = 1.310063
+ ags = 0.187311
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0018702
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.14095898
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 799951250.0
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.4509773e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.4407715
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.65 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.069866256e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.239906809e-8
+ k1 = 4.556237202e-01 lk1 = -6.484228401e-8
+ k2 = 2.007683582e-02 lk2 = 1.705422642e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.164179846e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.199470589e-8
+ nfactor = {2.378038919e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.167837078e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.443397737e-03 lu0 = 4.254027232e-9
+ ua = -7.572954228e-10 lua = 6.344807637e-16
+ ub = 8.922232633e-19 lub = -2.475144842e-25
+ uc = -7.084368051e-11 luc = -7.465141979e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.671623623e+05 lvsat = -8.547403617e-01 wvsat = 4.656612873e-16
+ a0 = 1.370094967e+00 la0 = -4.802116133e-7
+ ags = 1.321801322e-01 lags = 4.410064215e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.426888399e-04 lketa = -8.219334060e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.401119263e-01 lpclm = -7.931506930e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.387319811e-03 lpdiblc2 = 1.365168829e-08 wpdiblc2 = 8.673617380e-25 ppdiblc2 = 6.938893904e-30
+ pdiblcb = -2.488330300e-01 lpdiblcb = 7.496391204e-7
+ drout = 0.56
+ pscbe1 = 1.224636900e+09 lpscbe1 = -3.397173053e+3
+ pscbe2 = -1.698011262e-08 lpscbe2 = 1.792281353e-13 ppscbe2 = -5.293955920e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.446751046e+00 lbeta0 = 2.265262463e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.904539975e-10 lagidl = -1.962669803e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.670754974e+00 legidl = -6.281865390e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.063193317e-01 lkt1 = -2.755920237e-7
+ kt2 = -4.841666844e-02 lkt2 = -3.153153126e-8
+ at = -9.065933829e+04 lat = 7.252080717e-1
+ ute = -1.645263111e-01 lute = 2.580578176e-7
+ ua1 = 5.778773827e-10 lua1 = 9.957860376e-15
+ ub1 = 8.146409535e-19 lub1 = -1.224311373e-23 pub1 = -1.232595164e-44
+ uc1 = -1.163111597e-11 luc1 = 2.295664482e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.66 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063199473e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.736836213e-9
+ k1 = 4.427665361e-01 lk1 = -1.342299740e-8
+ k2 = 2.238297990e-02 lk2 = 7.831345119e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.585912374e-01 ldsub = -1.194145485e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.482687602e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.538498620e-8
+ nfactor = {9.059919706e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.719268760e-6
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394757071e-01 letab = 2.778517638e-7
+ u0 = 8.601632882e-03 lu0 = 3.621202956e-9
+ ua = -7.352853466e-10 lua = 5.464566366e-16 wua = -1.654361225e-30
+ ub = 8.528601283e-19 lub = -9.009087610e-26
+ uc = -7.556913799e-11 luc = 1.143321474e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.264314745e+00 la0 = -5.716847236e-8
+ ags = 1.560797535e-01 lags = 3.454255025e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.464757958e-03 lketa = -3.744375028e-08 wketa = 6.938893904e-24
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.488073345e-01 lpclm = 2.361946495e-06 ppclm = -1.332267630e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.621872386e-03 lpdiblc2 = -6.381398745e-09 wpdiblc2 = -6.938893904e-24
+ pdiblcb = -9.776424111e-02 lpdiblcb = 1.454750005e-7
+ drout = 0.56
+ pscbe1 = -4.171210305e+07 lpscbe1 = 1.667292191e+3
+ pscbe2 = 4.631193739e-08 lpscbe2 = -7.389354511e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.144527102e+01 lbeta0 = -9.335576356e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.690680066e-10 lagidl = -2.774355581e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815376811e-01 lkt1 = 2.522608815e-8
+ kt2 = -6.023855242e-02 lkt2 = 1.574731557e-8
+ at = 1.021557796e+05 lat = -4.591068088e-2
+ ute = -1.323451088e-01 lute = 1.293566616e-7
+ ua1 = 3.320607059e-09 lua1 = -1.011042424e-15
+ ub1 = -2.835183653e-18 lub1 = 2.353502076e-24
+ uc1 = 1.789645493e-11 luc1 = -9.513193603e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.67 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.080253346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.983204748e-8
+ k1 = 3.559763493e-01 lk1 = 1.600935854e-7
+ k2 = 5.664373486e-02 lk2 = -6.066498314e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.538016126e-01 ldsub = 1.029822606e-06 pdsub = 8.881784197e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.107617634e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.985602103e-10
+ nfactor = {2.269123695e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.992787282e-9
+ eta0 = -2.188386675e-01 leta0 = 4.385161211e-07 weta0 = 3.469446952e-24 peta0 = 1.804112415e-28
+ etab = 8.242798594e-01 letab = -1.648951009e-06 wetab = -1.058181320e-22 petab = 1.689620666e-27
+ u0 = 1.231769894e-02 lu0 = -3.808197859e-9
+ ua = -2.809317911e-10 lua = -3.619165246e-16
+ ub = 9.337272840e-19 lub = -2.517657501e-25
+ uc = -7.496753916e-11 luc = 1.023045924e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.949154737e+04 lvsat = -1.210264538e-2
+ a0 = 1.349266482e+00 la0 = -2.270095072e-7
+ ags = 1.615750419e-01 lags = 3.344389646e-7
+ a1 = 0.0
+ a2 = 6.001569927e-01 la2 = 3.995391301e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.083405179e-02 lketa = -2.858845418e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.592302506e-01 lpclm = 3.466122321e-7
+ pdiblc1 = 7.407420150e-01 lpdiblc1 = -7.012262346e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.203234000e-01 ldrout = 8.790300377e-7
+ pscbe1 = 7.981743154e+08 lpscbe1 = -1.186332945e+1
+ pscbe2 = 9.526279703e-09 lpscbe2 = -3.492672025e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.883960260e+00 lbeta0 = 1.782957602e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.471808281e-10 lagidl = 7.546826683e-16 pagidl = -4.135903063e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.587827164e-01 lkt1 = -2.026711633e-8
+ kt2 = -5.616202393e-02 lkt2 = 7.597254838e-9
+ at = 9.660944576e+04 lat = -3.482208970e-2
+ ute = 9.121531202e-01 lute = -1.958872090e-06 wute = -2.220446049e-22 pute = -2.220446049e-28
+ ua1 = 6.057818692e-09 lua1 = -6.483453838e-15 pua1 = 6.617444900e-36
+ ub1 = -4.209009179e-18 lub1 = 5.100143366e-24
+ uc1 = -1.262217768e-10 luc1 = 1.929986004e-16 wuc1 = -1.033975766e-31 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.68 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063768586e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.335940404e-8
+ k1 = 5.163411541e-01 lk1 = -1.533512796e-10
+ k2 = -5.168060475e-03 lk2 = 1.101380524e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.290252482e+00 ldsub = -5.130966086e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.913931266e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.895584058e-8
+ nfactor = {1.809580694e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.532124500e-7
+ eta0 = -4.960310000e-02 leta0 = 2.694049417e-7
+ etab = -1.649929909e+00 letab = 8.234402155e-7
+ u0 = 8.401454938e-03 lu0 = 1.051677069e-10
+ ua = -5.845179038e-10 lua = -5.855354765e-17
+ ub = 4.539112548e-19 lub = 2.276976143e-25
+ uc = -9.967858230e-11 luc = 3.492333976e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.063852456e+04 lvsat = 6.736520458e-3
+ a0 = 1.527093768e+00 la0 = -4.047060902e-7
+ ags = -2.563720022e-01 lags = 7.520788177e-7
+ a1 = 0.0
+ a2 = 1.009875667e+00 la2 = -9.878400712e-9
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.029268619e-02 lketa = -2.397005524e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.583204909e+00 lpclm = -7.765363053e-7
+ pdiblc1 = 6.695855342e-02 lpdiblc1 = -2.793800389e-8
+ pdiblc2 = 8.192914521e-04 lpdiblc2 = -3.890053229e-10
+ pdiblcb = -3.046280985e-02 lpdiblcb = 5.458794682e-9
+ drout = 1.0
+ pscbe1 = 7.726246557e+08 lpscbe1 = 1.366755128e+1
+ pscbe2 = 9.025583750e-09 lpscbe2 = 1.510607389e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.586477316e+00 lbeta0 = 1.080956896e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.230802340e-10 lagidl = -3.147917519e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.201462177e-01 lkt1 = -5.887521715e-8
+ kt2 = -6.442999755e-02 lkt2 = 1.585915150e-8
+ at = 8.839328001e+04 lat = -2.661196283e-2
+ ute = -1.896520674e+00 lute = 8.477373284e-07 pute = 1.776356839e-27
+ ua1 = -3.422902531e-09 lua1 = 2.990299055e-15 wua1 = -3.308722450e-30 pua1 = 2.481541838e-36
+ ub1 = 4.223470876e-18 lub1 = -3.326138816e-24 pub1 = 1.540743956e-45
+ uc1 = 3.287820583e-10 luc1 = -2.616708068e-16 wuc1 = 2.067951531e-31 puc1 = -2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.69 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.017357889e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.881673268e-10
+ k1 = 4.957720259e-01 lk1 = 1.011609452e-8
+ k2 = -1.259694042e-02 lk2 = 4.810360268e-09 wk2 = 6.938893904e-24 pk2 = -1.734723476e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.873419649e-01 ldsub = 2.745410829e-07 pdsub = -2.220446049e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.280419782e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.583516792e-10
+ nfactor = {2.822000291e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.225322040e-8
+ eta0 = 0.49
+ etab = -1.241930875e-03 letab = 3.080119933e-10
+ u0 = 1.000888135e-02 lu0 = -6.973640427e-10
+ ua = -1.854094572e-10 lua = -2.578144263e-16
+ ub = 2.788024247e-19 lub = 3.151233244e-25
+ uc = -5.941824113e-11 luc = 1.482276053e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.047205028e+04 lvsat = 1.680493524e-2
+ a0 = 8.395172334e-01 la0 = -6.142319168e-8
+ ags = 9.732161440e-01 lags = 1.381884919e-7
+ a1 = 0.0
+ a2 = 1.179620696e+00 la2 = -9.462615280e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.211104636e-02 lketa = 2.193294291e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.810947136e-01 lpclm = 3.040227459e-07 wpclm = 4.440892099e-22 ppclm = 1.387778781e-28
+ pdiblc1 = -3.856251289e-01 lpdiblc1 = 1.980211883e-07 wpdiblc1 = 1.387778781e-22 ppdiblc1 = -1.387778781e-29
+ pdiblc2 = -9.086226485e-03 lpdiblc2 = 4.556473090e-09 wpdiblc2 = 1.734723476e-24 ppdiblc2 = 1.544988096e-30
+ pdiblcb = 1.768499670e-01 lpdiblcb = -9.804521884e-08 wpdiblcb = -5.551115123e-23 ppdiblcb = 2.775557562e-29
+ drout = 1.509432333e+00 ldrout = -2.543417335e-7
+ pscbe1 = 8.000288649e+08 lpscbe1 = -1.441122781e-2
+ pscbe2 = 9.500903806e-09 lpscbe2 = -8.624992905e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.547070911e+00 lbeta0 = 1.021011347e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.848676046e-10 lagidl = -4.608102345e-17
+ bgidl = 7.403975816e+08 lbgidl = 1.296104014e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.586735669e-01 lkt1 = 1.028663983e-8
+ kt2 = -1.240616261e-02 lkt2 = -1.011452845e-8
+ at = -1.766680896e+03 lat = 1.840175005e-2
+ ute = 4.650627057e-01 lute = -3.313185975e-7
+ ua1 = 4.835890309e-09 lua1 = -1.133027153e-15
+ ub1 = -4.696559734e-18 lub1 = 1.127320267e-24
+ uc1 = -2.867396831e-10 luc1 = 4.563765543e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.70 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-4.324212251e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.456160701e-07 wvth0 = -4.698149683e-07 pvth0 = 1.171084281e-13
+ k1 = -3.689544462e+00 lk1 = 1.053369009e-06 wk1 = 3.647279892e-06 pk1 = -9.091392222e-13
+ k2 = 1.927008633e+00 lk2 = -4.786654230e-07 wk2 = -1.779151502e-06 pk2 = 4.434801992e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.543964640e+01 ldsub = -3.645646672e-06 wdsub = -1.731133297e-05 pdsub = 4.315109412e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {3.624761575e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.478538548e-07 wvoff = -4.128439965e-07 pvoff = 1.029075588e-13
+ nfactor = {-3.136350084e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.432954986e-06 wnfactor = 6.711219324e-06 pnfactor = -1.672872085e-12
+ eta0 = 6.457265625e+00 leta0 = -1.487430466e-06 weta0 = -6.598789180e-06 peta0 = 1.644847185e-12
+ etab = 6.272084162e-01 letab = -1.563426638e-07 wetab = -7.189836985e-07 petab = 1.792174716e-13
+ u0 = 2.110435616e-02 lu0 = -3.463077571e-09 wu0 = -5.524743947e-09 pu0 = 1.377125300e-15
+ ua = 1.590844829e-09 lua = -7.005724510e-16 wua = -5.619012267e-16 pua = 1.400623093e-22
+ ub = 3.700354112e-18 lub = -5.377497570e-25 wub = -3.844699063e-24 pub = 9.583489119e-31
+ uc = 1.803373179e-10 luc = -4.493990889e-17 wuc = -1.776702711e-16 puc = 4.428698012e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.234114606e+06 lvsat = -2.857136765e-01 wvsat = -1.394038306e+00 pvsat = 3.474849582e-7
+ a0 = 5.807526544e+00 la0 = -1.299774032e-06 wa0 = -6.924068830e-06 pa0 = 1.725928017e-12
+ ags = 2.238513771e+00 lags = -1.772059212e-7
+ a1 = 0.0
+ a2 = -5.278034159e-01 la2 = 3.309749185e-07 wa2 = 2.198657396e-06 pa2 = -5.480483359e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.759145120e-02 lketa = 8.544667402e-09 wketa = 9.092375064e-08 pketa = -2.266410870e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.802848148e-01 lpclm = 2.539678665e-07 wpclm = 1.035686253e-06 ppclm = -2.581603340e-13
+ pdiblc1 = 7.622584539e-01 lpdiblc1 = -8.810601300e-08 wpdiblc1 = -3.743552796e-07 ppdiblc1 = 9.331366878e-14
+ pdiblc2 = 5.624556379e-02 lpdiblc2 = -1.172845561e-08 wpdiblc2 = -5.612293728e-08 ppdiblc2 = 1.398948396e-14
+ pdiblcb = 1.720897528e+00 lpdiblcb = -4.829222341e-07 wpdiblcb = -2.464039307e-06 ppdiblcb = 6.141987578e-13
+ drout = -2.848517426e+00 ldrout = 8.319426132e-07 wdrout = 3.824438522e-06 pdrout = -9.532986681e-13
+ pscbe1 = 7.998969111e+08 lpscbe1 = 1.848022846e-2
+ pscbe2 = -4.502292578e-08 lpscbe2 = 1.350463245e-14 wpscbe2 = 6.943802332e-14 ppscbe2 = -1.730846888e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.752887417e+01 lbeta0 = -4.629398055e-06 wbeta0 = -2.216906880e-05 pbeta0 = 5.525972935e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.370563024e-08 lagidl = 8.426560422e-15 wagidl = 3.838581656e-14 pagidl = -9.568240564e-21
+ bgidl = 1.927151494e+09 lbgidl = -1.662058126e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.225139524e-01 lkt1 = -4.857968648e-08 wkt1 = -1.618340267e-07 pkt1 = 4.033955865e-14
+ kt2 = 1.599586990e-01 lkt2 = -5.307905568e-08 wkt2 = -2.733916157e-07 pkt2 = 6.814696109e-14
+ at = 6.412776943e+05 lat = -1.418867061e-01 wat = -5.912336440e-01 pat = 1.473738543e-7
+ ute = -1.706247212e+00 lute = 2.099129691e-07 wute = -8.442341724e-07 pute = 2.104380310e-13
+ ua1 = -5.016284362e-09 lua1 = 1.322775167e-15 wua1 = 6.364392822e-15 pua1 = -1.586420377e-21
+ ub1 = 1.044025482e-17 lub1 = -2.645757814e-24 wub1 = -1.375939867e-23 pub1 = 3.429736509e-30
+ uc1 = 1.265356699e-10 luc1 = -5.737742542e-17 wuc1 = -4.649491586e-16 puc1 = 1.158955520e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.71 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-2.409185905e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.285446341e-07 wvth0 = 1.681326201e-06 pvth0 = -2.939797054e-13
+ k1 = 8.264504785e+00 lk1 = -1.192899720e-06 wk1 = -9.242413337e-06 pk1 = 1.534441225e-12
+ k2 = -3.898477675e+00 lk2 = 6.192810041e-07 wk2 = 4.753468964e-06 pk2 = -7.965885870e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -3.654611728e+01 ldsub = 6.211616461e-06 wdsub = 4.747044296e-05 pdsub = -7.990076793e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.294960309e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.634216848e-07 wvoff = 1.232267098e-06 pvoff = -2.102112742e-13
+ nfactor = {2.635822000e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.219907293e-06 wnfactor = -3.027770246e-05 pnfactor = 5.428117389e-12
+ eta0 = -1.118018891e+01 leta0 = 1.833129027e-06 weta0 = 1.459096275e-05 peta0 = -2.357975865e-12
+ etab = -7.696916899e-01 letab = 1.029936991e-07 wetab = 9.557672527e-07 petab = -1.324820310e-13
+ u0 = 2.938473402e-02 lu0 = -5.416635373e-09 wu0 = -3.334306450e-08 pu0 = 6.967483080e-15
+ ua = 1.056505500e-08 lua = -2.528332267e-15 wua = -1.635116311e-14 pua = 3.252224135e-21
+ ub = -1.626889851e-17 lub = 3.330519900e-24 wub = 2.332936894e-23 pub = -4.284087714e-30
+ uc = 3.764778317e-10 luc = -8.769715361e-17 wuc = -5.053859233e-16 puc = 1.128059011e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.655775347e+06 lvsat = 4.506408690e-01 wvsat = 3.497828792e+00 pvsat = -5.796647575e-7
+ a0 = -1.387674807e+00 la0 = -1.086758636e-08 wa0 = 2.632508007e-06 pa0 = 1.397910675e-14
+ ags = 1.25
+ a1 = 0.0
+ a2 = 1.207243431e+01 la2 = -2.110623833e-06 wa2 = -1.469147300e-05 pa2 = 2.714920764e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.266105361e+00 lketa = -4.486680324e-07 wketa = -2.976054356e-06 pketa = 5.771270741e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.750110900e+00 lpclm = 5.469009810e-07 wpclm = 3.179946229e-06 ppclm = -7.034852947e-13
+ pdiblc1 = -1.085517800e+01 lpdiblc1 = 2.183634912e-06 wpdiblc1 = 1.445762470e-05 ppdiblc1 = -2.808835791e-12
+ pdiblc2 = -3.315423231e-01 lpdiblc2 = 6.326850493e-08 wpdiblc2 = 4.365740145e-07 ppdiblc2 = -8.138303711e-14
+ pdiblcb = -1.022365954e+01 lpdiblcb = 1.815579934e-06 wpdiblcb = 1.286139574e-05 ppdiblcb = -2.335402256e-12
+ drout = 2.495527201e+01 ldrout = -4.546073610e-06 wdrout = -3.128814199e-05 pdrout = 5.847669038e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 1.065860574e-07 lpscbe2 = -1.497023773e-14 wpscbe2 = -1.252286590e-13 ppscbe2 = 1.925639644e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -4.489186951e+01 lbeta0 = 9.145245637e-06 wbeta0 = 6.859418192e-05 pbeta0 = -1.176363921e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.744554069e-08 lagidl = -2.776169312e-15 wagidl = -3.318391178e-14 pagidl = 3.571019900e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.859125530e+00 lkt1 = 2.483964918e-07 wkt1 = 1.691172952e-06 pkt1 = -3.195153882e-13
+ kt2 = -2.552742778e+00 lkt2 = 4.742957241e-07 wkt2 = 3.215267763e-06 pkt2 = -6.100922814e-13
+ at = -1.462890967e+06 lat = 2.576326023e-01 wat = 1.919379412e+00 pat = -3.313959079e-7
+ ute = 1.047818369e+01 lute = -2.161557963e-06 wute = -1.383709446e-05 pute = 2.780437946e-12
+ ua1 = 2.727425018e-08 lua1 = -4.889285612e-15 wua1 = -3.452934794e-14 pua1 = 6.289146754e-21
+ ub1 = -4.248142011e-17 lub1 = 7.490013076e-24 wub1 = 5.446202574e-23 pub1 = -9.634493699e-30
+ uc1 = 4.061046702e-10 luc1 = -1.176882326e-16 wuc1 = -5.897684825e-16 puc1 = 1.513837858e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.72 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.109941926e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.824860809e-07 wvth0 = 1.776356839e-21
+ k1 = 4.276902357e-01 lk1 = 3.965345122e-7
+ k2 = 2.140283592e-02 lk2 = 1.611888913e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -2.094089633e-06 lcit = 2.418729035e-10 wcit = -8.470329473e-28 pcit = -4.065758147e-32
+ voff = {-2.660311031e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.622319741e-7
+ nfactor = {1.983358265e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.670632221e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.089193591e-02 lu0 = -3.833330944e-8
+ ua = -8.518531620e-10 lua = 3.477374642e-15
+ ub = 1.334168684e-18 lub = -9.457403913e-24
+ uc = -1.141341989e-10 luc = 8.471146658e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.011823641e+04 lvsat = 2.003761631e+0
+ a0 = 1.502482836e+00 la0 = -3.848255285e-6
+ ags = 9.478543007e-02 lags = 1.850443392e-6
+ a1 = 0.0
+ a2 = 1.012498438e+00 la2 = -4.249812576e-6
+ b0 = -1.621113085e-07 lb0 = 3.242107018e-12
+ b1 = 7.466570120e-10 lb1 = -1.493259145e-14
+ keta = 2.966889194e-02 lketa = -6.307586575e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.648858775e-02 lpclm = 3.148835631e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.516615195e-03 lpdiblc2 = -2.394546346e-8
+ pdiblcb = -2.424694755e-01 lpdiblcb = 1.746934707e-6
+ drout = 0.56
+ pscbe1 = 8.000121871e+08 lpscbe1 = -1.218696253e+0
+ pscbe2 = 1.121937296e-08 lpscbe2 = -1.158739448e-13
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.499908125e-11 lalpha0 = 2.499889751e-15
+ alpha1 = -2.499908125e-11 lalpha1 = 2.499889751e-15
+ beta0 = 3.593013473e+01 lbeta0 = -5.930091148e-04 pbeta0 = 9.094947018e-25
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.264033948e-09 lagidl = -3.637738745e-14 pagidl = 5.293955920e-35
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -9.635519618e-02 legidl = 1.963537530e-5
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.376196482e-01 lkt1 = -6.303472006e-8
+ kt2 = -6.009282515e-02 lkt2 = 1.546813783e-7
+ at = 8.873684778e+04 lat = -1.774671734e+0
+ ute = -7.065892282e-02 lute = -1.232098662e-6
+ ua1 = 2.157066468e-09 lua1 = -6.686597610e-15
+ ub1 = -1.357148067e-18 lub1 = 1.282471241e-23
+ uc1 = -3.504573888e-11 luc1 = 5.256700246e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.73 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.065816+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44751769
+ k2 = 0.02220881
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.22291792+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9820229+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0089752
+ ua = -6.7797804e-10
+ ub = 8.6128111e-19
+ uc = -7.1776909e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160310.0
+ a0 = 1.310063
+ ags = 0.187311
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0018702
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.14095898
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 799951250.0
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.4509773e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.4407715
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.74 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.069866256e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.239906809e-8
+ k1 = 4.556237202e-01 lk1 = -6.484228401e-8
+ k2 = 2.007683582e-02 lk2 = 1.705422642e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.164179846e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.199470589e-8
+ nfactor = {2.378038919e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.167837078e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.443397737e-03 lu0 = 4.254027232e-9
+ ua = -7.572954228e-10 lua = 6.344807637e-16
+ ub = 8.922232633e-19 lub = -2.475144842e-25
+ uc = -7.084368051e-11 luc = -7.465141979e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.671623623e+05 lvsat = -8.547403617e-1
+ a0 = 1.370094967e+00 la0 = -4.802116133e-7
+ ags = 1.321801322e-01 lags = 4.410064215e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.426888399e-04 lketa = -8.219334060e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.401119263e-01 lpclm = -7.931506930e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.387319811e-03 lpdiblc2 = 1.365168829e-08 wpdiblc2 = -8.673617380e-25 ppdiblc2 = 6.938893904e-30
+ pdiblcb = -2.488330300e-01 lpdiblcb = 7.496391204e-7
+ drout = 0.56
+ pscbe1 = 1.224636900e+09 lpscbe1 = -3.397173053e+3
+ pscbe2 = -1.698011262e-08 lpscbe2 = 1.792281353e-13 wpscbe2 = -1.323488980e-29
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.446751046e+00 lbeta0 = 2.265262463e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.904539975e-10 lagidl = -1.962669803e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.670754974e+00 legidl = -6.281865390e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.063193317e-01 lkt1 = -2.755920237e-7
+ kt2 = -4.841666844e-02 lkt2 = -3.153153126e-8
+ at = -9.065933829e+04 lat = 7.252080717e-1
+ ute = -1.645263111e-01 lute = 2.580578176e-7
+ ua1 = 5.778773827e-10 lua1 = 9.957860376e-15
+ ub1 = 8.146409535e-19 lub1 = -1.224311373e-23 pub1 = -1.232595164e-44
+ uc1 = -1.163111597e-11 luc1 = 2.295664482e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.75 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063199473e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.736836213e-9
+ k1 = 4.427665361e-01 lk1 = -1.342299740e-8
+ k2 = 2.238297990e-02 lk2 = 7.831345119e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.585912374e-01 ldsub = -1.194145485e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.482687602e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.538498620e-8
+ nfactor = {9.059919706e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.719268760e-6
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394757071e-01 letab = 2.778517638e-7
+ u0 = 8.601632882e-03 lu0 = 3.621202956e-9
+ ua = -7.352853466e-10 lua = 5.464566366e-16
+ ub = 8.528601283e-19 lub = -9.009087610e-26
+ uc = -7.556913799e-11 luc = 1.143321474e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.264314745e+00 la0 = -5.716847236e-8
+ ags = 1.560797535e-01 lags = 3.454255025e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.464757958e-03 lketa = -3.744375028e-08 wketa = 6.938893904e-24 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.488073345e-01 lpclm = 2.361946495e-06 wpclm = 1.110223025e-22 ppclm = -1.110223025e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.621872386e-03 lpdiblc2 = -6.381398745e-9
+ pdiblcb = -9.776424111e-02 lpdiblcb = 1.454750005e-7
+ drout = 0.56
+ pscbe1 = -4.171210305e+07 lpscbe1 = 1.667292191e+3
+ pscbe2 = 4.631193739e-08 lpscbe2 = -7.389354511e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.144527102e+01 lbeta0 = -9.335576356e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.690680066e-10 lagidl = -2.774355581e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815376811e-01 lkt1 = 2.522608815e-8
+ kt2 = -6.023855242e-02 lkt2 = 1.574731557e-8
+ at = 1.021557796e+05 lat = -4.591068088e-2
+ ute = -1.323451088e-01 lute = 1.293566616e-7
+ ua1 = 3.320607059e-09 lua1 = -1.011042424e-15
+ ub1 = -2.835183653e-18 lub1 = 2.353502076e-24
+ uc1 = 1.789645493e-11 luc1 = -9.513193603e-17 puc1 = 7.754818243e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.76 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.080253346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.983204748e-8
+ k1 = 3.559763493e-01 lk1 = 1.600935854e-7
+ k2 = 5.664373486e-02 lk2 = -6.066498314e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.538016126e-01 ldsub = 1.029822606e-06 pdsub = 8.881784197e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.107617634e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.985602103e-10
+ nfactor = {2.269123695e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.992787282e-9
+ eta0 = -2.188386675e-01 leta0 = 4.385161211e-07 weta0 = 2.775557562e-23 peta0 = 1.387778781e-29
+ etab = 8.242798594e-01 letab = -1.648951009e-06 wetab = -2.428612866e-23 petab = -1.179611964e-27
+ u0 = 1.231769894e-02 lu0 = -3.808197859e-9
+ ua = -2.809317911e-10 lua = -3.619165246e-16
+ ub = 9.337272840e-19 lub = -2.517657501e-25
+ uc = -7.496753916e-11 luc = 1.023045924e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.949154737e+04 lvsat = -1.210264538e-2
+ a0 = 1.349266482e+00 la0 = -2.270095072e-7
+ ags = 1.615750419e-01 lags = 3.344389646e-7
+ a1 = 0.0
+ a2 = 6.001569927e-01 la2 = 3.995391301e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.083405178e-02 lketa = -2.858845418e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.592302506e-01 lpclm = 3.466122321e-7
+ pdiblc1 = 7.407420150e-01 lpdiblc1 = -7.012262346e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.203234000e-01 ldrout = 8.790300377e-7
+ pscbe1 = 7.981743154e+08 lpscbe1 = -1.186332945e+1
+ pscbe2 = 9.526279703e-09 lpscbe2 = -3.492672025e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.883960260e+00 lbeta0 = 1.782957602e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.471808281e-10 lagidl = 7.546826683e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.587827164e-01 lkt1 = -2.026711633e-8
+ kt2 = -5.616202393e-02 lkt2 = 7.597254838e-9
+ at = 9.660944576e+04 lat = -3.482208970e-2
+ ute = 9.121531202e-01 lute = -1.958872090e-06 wute = 6.661338148e-22 pute = -6.661338148e-28
+ ua1 = 6.057818692e-09 lua1 = -6.483453838e-15
+ ub1 = -4.209009179e-18 lub1 = 5.100143366e-24 wub1 = -6.162975822e-39
+ uc1 = -1.262217768e-10 luc1 = 1.929986004e-16 wuc1 = -1.033975766e-31 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.77 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063768586e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.335940404e-8
+ k1 = 5.163411541e-01 lk1 = -1.533512796e-10
+ k2 = -5.168060475e-03 lk2 = 1.101380524e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.290252482e+00 ldsub = -5.130966086e-07 wdsub = -1.776356839e-21
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.913931266e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.895584058e-8
+ nfactor = {1.809580694e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.532124500e-7
+ eta0 = -4.960310000e-02 leta0 = 2.694049417e-7
+ etab = -1.649929909e+00 letab = 8.234402155e-7
+ u0 = 8.401454938e-03 lu0 = 1.051677069e-10
+ ua = -5.845179038e-10 lua = -5.855354765e-17
+ ub = 4.539112548e-19 lub = 2.276976143e-25
+ uc = -9.967858230e-11 luc = 3.492333976e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.063852456e+04 lvsat = 6.736520458e-3
+ a0 = 1.527093768e+00 la0 = -4.047060902e-7
+ ags = -2.563720022e-01 lags = 7.520788177e-7
+ a1 = 0.0
+ a2 = 1.009875667e+00 la2 = -9.878400712e-9
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.029268619e-02 lketa = -2.397005524e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.583204909e+00 lpclm = -7.765363053e-7
+ pdiblc1 = 6.695855342e-02 lpdiblc1 = -2.793800389e-8
+ pdiblc2 = 8.192914521e-04 lpdiblc2 = -3.890053229e-10
+ pdiblcb = -3.046280985e-02 lpdiblcb = 5.458794682e-9
+ drout = 1.0
+ pscbe1 = 7.726246557e+08 lpscbe1 = 1.366755128e+1
+ pscbe2 = 9.025583750e-09 lpscbe2 = 1.510607389e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.586477316e+00 lbeta0 = 1.080956896e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.230802340e-10 lagidl = -3.147917519e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.201462177e-01 lkt1 = -5.887521715e-8
+ kt2 = -6.442999755e-02 lkt2 = 1.585915150e-8
+ at = 8.839328001e+04 lat = -2.661196283e-2
+ ute = -1.896520674e+00 lute = 8.477373284e-7
+ ua1 = -3.422902531e-09 lua1 = 2.990299055e-15 pua1 = -8.271806126e-37
+ ub1 = 4.223470876e-18 lub1 = -3.326138816e-24 pub1 = 1.540743956e-45
+ uc1 = 3.287820583e-10 luc1 = -2.616708068e-16 wuc1 = -2.067951531e-31 puc1 = -2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.78 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.017357889e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.881673268e-10
+ k1 = 4.957720259e-01 lk1 = 1.011609452e-8
+ k2 = -1.259694042e-02 lk2 = 4.810360268e-09 wk2 = 6.938893904e-24 pk2 = -1.734723476e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.873419649e-01 ldsub = 2.745410829e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.280419782e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.583516792e-10
+ nfactor = {2.822000291e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.225322040e-8
+ eta0 = 0.49
+ etab = -1.241930875e-03 letab = 3.080119933e-10
+ u0 = 1.000888135e-02 lu0 = -6.973640427e-10
+ ua = -1.854094572e-10 lua = -2.578144263e-16
+ ub = 2.788024247e-19 lub = 3.151233244e-25
+ uc = -5.941824113e-11 luc = 1.482276053e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.047205028e+04 lvsat = 1.680493524e-2
+ a0 = 8.395172334e-01 la0 = -6.142319168e-08 wa0 = 1.776356839e-21
+ ags = 9.732161440e-01 lags = 1.381884919e-7
+ a1 = 0.0
+ a2 = 1.179620696e+00 la2 = -9.462615280e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.211104636e-02 lketa = 2.193294291e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.810947136e-01 lpclm = 3.040227459e-07 wpclm = 3.330669074e-22 ppclm = 5.551115123e-29
+ pdiblc1 = -3.856251289e-01 lpdiblc1 = 1.980211883e-07 wpdiblc1 = 1.942890293e-22 ppdiblc1 = 6.245004514e-29
+ pdiblc2 = -9.086226485e-03 lpdiblc2 = 4.556473090e-09 ppdiblc2 = -2.927345866e-30
+ pdiblcb = 1.768499670e-01 lpdiblcb = -9.804521884e-08 wpdiblcb = 5.551115123e-23 ppdiblcb = 4.163336342e-29
+ drout = 1.509432333e+00 ldrout = -2.543417335e-7
+ pscbe1 = 8.000288649e+08 lpscbe1 = -1.441122781e-2
+ pscbe2 = 9.500903806e-09 lpscbe2 = -8.624992905e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.547070911e+00 lbeta0 = 1.021011347e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.848676046e-10 lagidl = -4.608102345e-17
+ bgidl = 7.403975816e+08 lbgidl = 1.296104014e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.586735669e-01 lkt1 = 1.028663983e-8
+ kt2 = -1.240616261e-02 lkt2 = -1.011452845e-8
+ at = -1.766680896e+03 lat = 1.840175005e-2
+ ute = 4.650627057e-01 lute = -3.313185975e-07 wute = -4.440892099e-22 pute = 1.110223025e-28
+ ua1 = 4.835890309e-09 lua1 = -1.133027153e-15
+ ub1 = -4.696559734e-18 lub1 = 1.127320267e-24 pub1 = -1.540743956e-45
+ uc1 = -2.867396831e-10 luc1 = 4.563765543e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.79 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.422703484e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.345502839e-8
+ k1 = -5.077929917e-01 lk1 = 2.602697286e-7
+ k2 = 3.749429630e-01 lk2 = -9.178977375e-08 wk2 = 8.326672685e-23 pk2 = 6.938893904e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.378826863e-01 ldsub = 1.186944602e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {2.326393325e-03+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.808112382e-8
+ nfactor = {2.718268313e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.639646891e-8
+ eta0 = 7.007271087e-01 leta0 = -5.252689275e-8
+ etab = -6.25e-6
+ u0 = 1.628477480e-02 lu0 = -2.261724623e-9
+ ua = 1.100663075e-09 lua = -5.783872961e-16
+ ub = 3.463814915e-19 lub = 2.982782283e-25
+ uc = 2.534437437e-11 luc = -6.305592823e-18 wuc = -1.494418099e-32 puc = 4.038967835e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.800738114e+04 lvsat = 1.741929099e-2
+ a0 = -2.327738550e-01 la0 = 2.058614465e-7
+ ags = 2.238513771e+00 lags = -1.772059212e-7
+ a1 = 0.0
+ a2 = 1.390223610e+00 la2 = -1.471220882e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.172705079e-02 lketa = -1.122665899e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.232093940e-01 lpclm = 2.875838254e-8
+ pdiblc1 = 4.356848163e-01 lpdiblc1 = -6.702635233e-9
+ pdiblc2 = 7.285998437e-03 lpdiblc2 = 4.754504447e-10
+ pdiblcb = -4.286388172e-01 lpdiblcb = 5.288194294e-8
+ drout = 4.877806509e-01 ldrout = 3.202728919e-10
+ pscbe1 = 7.998969111e+08 lpscbe1 = 1.848022846e-2
+ pscbe2 = 1.555222594e-08 lpscbe2 = -1.594632741e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.189402196e+00 lbeta0 = 1.912554271e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.192700175e-10 lagidl = 7.958284090e-17
+ bgidl = 1.927151494e+09 lbgidl = -1.662058126e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.636919446e-01 lkt1 = -1.338895424e-8
+ kt2 = -7.853798926e-02 lkt2 = 6.369821319e-9
+ at = 1.255074293e+05 lat = -1.332323102e-2
+ ute = -2.442725738e+00 lute = 3.934912890e-7
+ ua1 = 5.357754802e-10 lua1 = -6.115902980e-17
+ ub1 = -1.562933375e-18 lub1 = 3.462168921e-25 wub1 = -1.540743956e-39
+ uc1 = -2.790687019e-10 luc1 = 4.372554830e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.80 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-9.424588082e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.791245342e-08 wvth0 = -6.701769024e-13 pvth0 = 1.315322695e-19
+ k1 = 2.017663331e-01 lk1 = 1.456898817e-07 wk1 = 5.037250830e-13 pk1 = -9.886360353e-20
+ k2 = 2.482719274e-01 lk2 = -7.563326083e-08 wk2 = 1.328939092e-13 pk2 = -2.608242289e-20
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.865334068e+00 ldsub = -7.586297909e-07 wdsub = -6.542595372e-13 pdsub = 1.284082476e-19
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.199761962e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.995883628e-08 wvoff = -8.996905621e-14 pvoff = 1.765777746e-20
+ nfactor = {-5.496894413e-02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.153897201e-07 wnfactor = 5.298900163e-11 pnfactor = -1.039988641e-17
+ eta0 = 1.548433626e+00 leta0 = -2.238832255e-07 weta0 = -1.000761765e-11 peta0 = 1.964145077e-18
+ etab = 6.408315235e-02 letab = -1.257850655e-08 wetab = 1.145733678e-12 petab = -2.248674204e-19
+ u0 = 2.974684976e-04 lu0 = 6.615409171e-10 wu0 = 1.701528973e-14 pu0 = -3.339505845e-21
+ ua = -3.699095870e-09 lua = 3.087879580e-16 wua = 4.199882082e-21 pua = -8.242898545e-28
+ ub = 4.082756185e-18 lub = -4.067551273e-25 wub = 2.294101047e-29 pub = -4.502517417e-36
+ uc = -6.440236335e-11 luc = 1.071058073e-17 wuc = 3.348320459e-22 puc = -6.571581150e-29
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.956004339e+05 lvsat = -5.503710899e-02 wvsat = 1.181412945e-07 pvsat = -2.318700124e-14
+ a0 = 9.088172489e-01 la0 = 1.329253988e-09 wa0 = 1.160526038e-11 pa0 = -2.277706429e-18
+ ags = 1.25
+ a1 = 0.0
+ a2 = -7.438583539e-01 la2 = 2.577716746e-07 wa2 = -2.918594348e-12 pa2 = 5.728179193e-19
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.300942480e-01 lketa = 5.479625536e-08 wketa = 4.103245583e-13 pketa = -8.053234946e-20
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.023954717e+00 lpclm = -6.679319280e-08 wpclm = 1.523035351e-12 ppclm = -2.989185344e-19
+ pdiblc1 = 1.757129295e+00 lpdiblc1 = -2.666915579e-07 wpdiblc1 = -1.449823240e-11 ppdiblc1 = 2.845495582e-18
+ pdiblc2 = 4.930844220e-02 lpdiblc2 = -7.726996719e-09 wpdiblc2 = 2.120923784e-13 ppdiblc2 = -4.162631065e-20
+ pdiblcb = 9.961049512e-01 lpdiblcb = -2.217305096e-07 wpdiblcb = 4.507615183e-11 ppdiblcb = -8.846870939e-18
+ drout = -2.339378494e+00 ldrout = 5.552230345e-07 wdrout = 4.341911234e-11 pdrout = -8.521652083e-18
+ pscbe1 = 800000000.0
+ pscbe2 = -2.658580395e-09 lpscbe2 = 1.828289472e-15 wpscbe2 = -2.197075702e-19 ppscbe2 = 4.312090626e-26
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.494712325e+01 lbeta0 = -1.116911624e-06 wbeta0 = 2.645067468e-11 pbeta0 = -5.191341671e-18
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.503194015e-09 lagidl = 3.391191583e-16 wagidl = 3.701981390e-19 pagidl = -7.265693775e-26
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.838099919e-01 lkt1 = -3.033668264e-08 wkt1 = 1.047059378e-12 pkt1 = -2.055011095e-19
+ kt2 = 2.521358021e-01 lkt2 = -5.792580953e-08 wkt2 = 1.787345545e-12 pkt2 = -3.507933735e-19
+ at = 2.115048933e+05 lat = -3.146498760e-02 wat = -6.549507030e-07 pat = 1.285438997e-13
+ ute = -1.592779878e+00 lute = 2.639921023e-07 wute = -4.076300348e-12 pute = 8.000350875e-19
+ ua1 = -2.847843263e-09 lua1 = 5.971270897e-16 wua1 = -3.076034822e-20 pua1 = 6.037179742e-27
+ ub1 = 5.029196934e-18 lub1 = -9.147552355e-25 wub1 = 3.529427768e-29 pub1 = -6.927031409e-36
+ uc1 = -1.083895978e-10 luc1 = 1.437378086e-17 wuc1 = 2.470778633e-21 puc1 = -4.849273685e-28
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.81 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.109941926e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.824860809e-7
+ k1 = 4.276902357e-01 lk1 = 3.965345122e-7
+ k2 = 2.140283592e-02 lk2 = 1.611888913e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -2.094089633e-06 lcit = 2.418729035e-10 pcit = -1.355252716e-31
+ voff = {-2.660311031e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.622319741e-7
+ nfactor = {1.983358265e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.670632221e-08 wnfactor = -7.105427358e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.089193591e-02 lu0 = -3.833330944e-8
+ ua = -8.518531620e-10 lua = 3.477374642e-15
+ ub = 1.334168684e-18 lub = -9.457403913e-24
+ uc = -1.141341989e-10 luc = 8.471146658e-16 wuc = -4.135903063e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.011823641e+04 lvsat = 2.003761631e+0
+ a0 = 1.502482836e+00 la0 = -3.848255285e-6
+ ags = 9.478543007e-02 lags = 1.850443392e-6
+ a1 = 0.0
+ a2 = 1.012498438e+00 la2 = -4.249812576e-6
+ b0 = -1.621113085e-07 lb0 = 3.242107018e-12
+ b1 = 7.466570120e-10 lb1 = -1.493259145e-14
+ keta = 2.966889194e-02 lketa = -6.307586575e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.648858775e-02 lpclm = 3.148835631e-06 ppclm = 2.664535259e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.516615195e-03 lpdiblc2 = -2.394546346e-8
+ pdiblcb = -2.424694755e-01 lpdiblcb = 1.746934707e-6
+ drout = 0.56
+ pscbe1 = 8.000121871e+08 lpscbe1 = -1.218696253e+0
+ pscbe2 = 1.121937296e-08 lpscbe2 = -1.158739448e-13
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.499908125e-11 lalpha0 = 2.499889751e-15
+ alpha1 = -2.499908125e-11 lalpha1 = 2.499889751e-15
+ beta0 = 3.593013473e+01 lbeta0 = -5.930091148e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.264033948e-09 lagidl = -3.637738745e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -9.635519618e-02 legidl = 1.963537530e-05 pegidl = -1.421085472e-26
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.376196482e-01 lkt1 = -6.303472006e-8
+ kt2 = -6.009282515e-02 lkt2 = 1.546813783e-7
+ at = 8.873684778e+04 lat = -1.774671734e+0
+ ute = -7.065892282e-02 lute = -1.232098662e-6
+ ua1 = 2.157066468e-09 lua1 = -6.686597610e-15
+ ub1 = -1.357148067e-18 lub1 = 1.282471241e-23
+ uc1 = -3.504573888e-11 luc1 = 5.256700246e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.82 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.065816+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44751769
+ k2 = 0.02220881
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.22291792+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9820229+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0089752
+ ua = -6.7797804e-10
+ ub = 8.6128111e-19
+ uc = -7.1776909e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160310.0
+ a0 = 1.310063
+ ags = 0.187311
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0018702
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.14095898
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 799951250.0
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.4509773e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.4407715
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.83 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.069866256e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.239906809e-8
+ k1 = 4.556237202e-01 lk1 = -6.484228401e-8
+ k2 = 2.007683582e-02 lk2 = 1.705422642e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.164179846e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.199470589e-8
+ nfactor = {2.378038919e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.167837078e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.443397737e-03 lu0 = 4.254027232e-9
+ ua = -7.572954228e-10 lua = 6.344807637e-16
+ ub = 8.922232633e-19 lub = -2.475144842e-25
+ uc = -7.084368051e-11 luc = -7.465141979e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.671623623e+05 lvsat = -8.547403617e-1
+ a0 = 1.370094967e+00 la0 = -4.802116133e-7
+ ags = 1.321801322e-01 lags = 4.410064215e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.426888399e-04 lketa = -8.219334060e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.401119263e-01 lpclm = -7.931506930e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.387319811e-03 lpdiblc2 = 1.365168829e-08 wpdiblc2 = -1.734723476e-24 ppdiblc2 = -6.938893904e-30
+ pdiblcb = -2.488330300e-01 lpdiblcb = 7.496391204e-7
+ drout = 0.56
+ pscbe1 = 1.224636900e+09 lpscbe1 = -3.397173053e+03 wpscbe1 = -3.814697266e-12
+ pscbe2 = -1.698011262e-08 lpscbe2 = 1.792281353e-13 ppscbe2 = -1.058791184e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.446751046e+00 lbeta0 = 2.265262463e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.904539975e-10 lagidl = -1.962669803e-15 pagidl = -6.617444900e-36
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.670754974e+00 legidl = -6.281865390e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.063193317e-01 lkt1 = -2.755920237e-7
+ kt2 = -4.841666844e-02 lkt2 = -3.153153126e-8
+ at = -9.065933828e+04 lat = 7.252080717e-1
+ ute = -1.645263111e-01 lute = 2.580578176e-7
+ ua1 = 5.778773827e-10 lua1 = 9.957860376e-15
+ ub1 = 8.146409535e-19 lub1 = -1.224311373e-23 pub1 = 1.232595164e-44
+ uc1 = -1.163111597e-11 luc1 = 2.295664482e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.84 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063199473e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.736836213e-9
+ k1 = 4.427665361e-01 lk1 = -1.342299740e-8
+ k2 = 2.238297990e-02 lk2 = 7.831345119e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.585912374e-01 ldsub = -1.194145485e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.482687602e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.538498620e-8
+ nfactor = {9.059919706e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.719268760e-6
+ eta0 = 1.594707837e-01 leta0 = -3.178247240e-7
+ etab = -1.394757071e-01 letab = 2.778517638e-7
+ u0 = 8.601632881e-03 lu0 = 3.621202956e-9
+ ua = -7.352853466e-10 lua = 5.464566366e-16
+ ub = 8.528601283e-19 lub = -9.009087610e-26
+ uc = -7.556913799e-11 luc = 1.143321474e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.264314745e+00 la0 = -5.716847236e-8
+ ags = 1.560797535e-01 lags = 3.454255025e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.464757958e-03 lketa = -3.744375028e-08 pketa = 5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.488073345e-01 lpclm = 2.361946495e-06 wpclm = 8.881784197e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.621872386e-03 lpdiblc2 = -6.381398745e-9
+ pdiblcb = -9.776424111e-02 lpdiblcb = 1.454750005e-7
+ drout = 0.56
+ pscbe1 = -4.171210305e+07 lpscbe1 = 1.667292191e+3
+ pscbe2 = 4.631193739e-08 lpscbe2 = -7.389354511e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.144527102e+01 lbeta0 = -9.335576356e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.690680066e-10 lagidl = -2.774355581e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815376811e-01 lkt1 = 2.522608815e-8
+ kt2 = -6.023855242e-02 lkt2 = 1.574731557e-8
+ at = 1.021557796e+05 lat = -4.591068088e-2
+ ute = -1.323451088e-01 lute = 1.293566616e-7
+ ua1 = 3.320607059e-09 lua1 = -1.011042424e-15
+ ub1 = -2.835183653e-18 lub1 = 2.353502076e-24
+ uc1 = 1.789645493e-11 luc1 = -9.513193603e-17 wuc1 = -2.584939414e-32 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.85 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.080253346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.983204748e-8
+ k1 = 3.559763493e-01 lk1 = 1.600935854e-7
+ k2 = 5.664373486e-02 lk2 = -6.066498314e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.538016126e-01 ldsub = 1.029822606e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.107617634e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.985602103e-10
+ nfactor = {2.269123695e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.992787282e-9
+ eta0 = -2.188386675e-01 leta0 = 4.385161211e-07 weta0 = -1.075528555e-22 peta0 = 9.367506770e-29
+ etab = 8.242798594e-01 letab = -1.648951009e-06 wetab = -5.065392550e-22 petab = 8.743006319e-28
+ u0 = 1.231769894e-02 lu0 = -3.808197859e-9
+ ua = -2.809317911e-10 lua = -3.619165246e-16
+ ub = 9.337272840e-19 lub = -2.517657501e-25
+ uc = -7.496753916e-11 luc = 1.023045924e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.949154737e+04 lvsat = -1.210264538e-2
+ a0 = 1.349266482e+00 la0 = -2.270095072e-7
+ ags = 1.615750419e-01 lags = 3.344389646e-7
+ a1 = 0.0
+ a2 = 6.001569926e-01 la2 = 3.995391301e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.083405179e-02 lketa = -2.858845418e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.592302506e-01 lpclm = 3.466122321e-7
+ pdiblc1 = 7.407420150e-01 lpdiblc1 = -7.012262346e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.203234000e-01 ldrout = 8.790300377e-7
+ pscbe1 = 7.981743154e+08 lpscbe1 = -1.186332945e+1
+ pscbe2 = 9.526279703e-09 lpscbe2 = -3.492672025e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.883960260e+00 lbeta0 = 1.782957602e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.471808281e-10 lagidl = 7.546826683e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.587827164e-01 lkt1 = -2.026711633e-8
+ kt2 = -5.616202393e-02 lkt2 = 7.597254838e-9
+ at = 9.660944576e+04 lat = -3.482208970e-2
+ ute = 9.121531202e-01 lute = -1.958872090e-06 wute = 4.440892099e-22 pute = -2.220446049e-27
+ ua1 = 6.057818692e-09 lua1 = -6.483453838e-15
+ ub1 = -4.209009179e-18 lub1 = 5.100143366e-24 wub1 = -6.162975822e-39 pub1 = -6.162975822e-45
+ uc1 = -1.262217768e-10 luc1 = 1.929986004e-16 wuc1 = -2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.86 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063768586e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.335940404e-8
+ k1 = 5.163411541e-01 lk1 = -1.533512796e-10
+ k2 = -5.168060475e-03 lk2 = 1.101380524e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.290252482e+00 ldsub = -5.130966086e-07 pdsub = 1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.913931266e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.895584058e-8
+ nfactor = {1.809580694e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.532124500e-7
+ eta0 = -4.960310000e-02 leta0 = 2.694049417e-7
+ etab = -1.649929909e+00 letab = 8.234402155e-7
+ u0 = 8.401454938e-03 lu0 = 1.051677069e-10
+ ua = -5.845179038e-10 lua = -5.855354765e-17
+ ub = 4.539112548e-19 lub = 2.276976143e-25
+ uc = -9.967858230e-11 luc = 3.492333976e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.063852456e+04 lvsat = 6.736520458e-3
+ a0 = 1.527093768e+00 la0 = -4.047060902e-7
+ ags = -2.563720022e-01 lags = 7.520788177e-7
+ a1 = 0.0
+ a2 = 1.009875667e+00 la2 = -9.878400712e-9
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.029268619e-02 lketa = -2.397005524e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.583204909e+00 lpclm = -7.765363053e-7
+ pdiblc1 = 6.695855342e-02 lpdiblc1 = -2.793800389e-08 wpdiblc1 = 2.220446049e-22
+ pdiblc2 = 8.192914521e-04 lpdiblc2 = -3.890053229e-10
+ pdiblcb = -3.046280985e-02 lpdiblcb = 5.458794682e-9
+ drout = 1.0
+ pscbe1 = 7.726246557e+08 lpscbe1 = 1.366755128e+1
+ pscbe2 = 9.025583750e-09 lpscbe2 = 1.510607389e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.586477316e+00 lbeta0 = 1.080956896e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.230802340e-10 lagidl = -3.147917519e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.201462177e-01 lkt1 = -5.887521715e-8
+ kt2 = -6.442999755e-02 lkt2 = 1.585915150e-08 wkt2 = 2.220446049e-22
+ at = 8.839328001e+04 lat = -2.661196283e-02 wat = 2.328306437e-16
+ ute = -1.896520674e+00 lute = 8.477373284e-7
+ ua1 = -3.422902531e-09 lua1 = 2.990299055e-15 wua1 = 1.654361225e-30 pua1 = 1.654361225e-36
+ ub1 = 4.223470876e-18 lub1 = -3.326138816e-24 pub1 = -3.081487911e-45
+ uc1 = 3.287820583e-10 luc1 = -2.616708068e-16 wuc1 = 4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.87 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.017357889e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.881673268e-10
+ k1 = 4.957720259e-01 lk1 = 1.011609452e-8
+ k2 = -1.259694042e-02 lk2 = 4.810360268e-09 wk2 = -1.387778781e-23 pk2 = 3.469446952e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.873419649e-01 ldsub = 2.745410829e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.280419782e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.583516792e-10
+ nfactor = {2.822000291e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.225322040e-8
+ eta0 = 0.49
+ etab = -1.241930875e-03 letab = 3.080119933e-10
+ u0 = 1.000888135e-02 lu0 = -6.973640427e-10
+ ua = -1.854094572e-10 lua = -2.578144263e-16
+ ub = 2.788024247e-19 lub = 3.151233244e-25
+ uc = -5.941824113e-11 luc = 1.482276053e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.047205028e+04 lvsat = 1.680493524e-2
+ a0 = 8.395172334e-01 la0 = -6.142319168e-8
+ ags = 9.732161440e-01 lags = 1.381884919e-7
+ a1 = 0.0
+ a2 = 1.179620696e+00 la2 = -9.462615280e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.211104636e-02 lketa = 2.193294291e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.810947136e-01 lpclm = 3.040227459e-07 wpclm = -1.110223025e-22 ppclm = -2.498001805e-28
+ pdiblc1 = -3.856251289e-01 lpdiblc1 = 1.980211883e-07 wpdiblc1 = -3.330669074e-22 ppdiblc1 = 1.387778781e-28
+ pdiblc2 = -9.086226485e-03 lpdiblc2 = 4.556473090e-09 wpdiblc2 = 1.149254303e-23 ppdiblc2 = 2.059984128e-30
+ pdiblcb = 1.768499670e-01 lpdiblcb = -9.804521884e-08 wpdiblcb = -1.110223025e-22 ppdiblcb = 2.775557562e-29
+ drout = 1.509432333e+00 ldrout = -2.543417335e-7
+ pscbe1 = 8.000288649e+08 lpscbe1 = -1.441122781e-2
+ pscbe2 = 9.500903806e-09 lpscbe2 = -8.624992905e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.547070911e+00 lbeta0 = 1.021011347e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.848676046e-10 lagidl = -4.608102345e-17
+ bgidl = 7.403975816e+08 lbgidl = 1.296104014e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.586735669e-01 lkt1 = 1.028663983e-8
+ kt2 = -1.240616261e-02 lkt2 = -1.011452845e-8
+ at = -1.766680896e+03 lat = 1.840175005e-2
+ ute = 4.650627057e-01 lute = -3.313185975e-07 pute = 2.220446049e-28
+ ua1 = 4.835890309e-09 lua1 = -1.133027153e-15
+ ub1 = -4.696559734e-18 lub1 = 1.127320267e-24 wub1 = 1.232595164e-38
+ uc1 = -2.867396831e-10 luc1 = 4.563765543e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.88 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.422703484e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.345502839e-8
+ k1 = -5.077929916e-01 lk1 = 2.602697286e-7
+ k2 = 3.749429630e-01 lk2 = -9.178977375e-08 wk2 = 1.665334537e-22 pk2 = -1.387778781e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.378826863e-01 ldsub = 1.186944602e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {2.326393325e-03+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.808112382e-8
+ nfactor = {2.718268313e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.639646891e-8
+ eta0 = 7.007271087e-01 leta0 = -5.252689275e-8
+ etab = -6.25e-6
+ u0 = 1.628477480e-02 lu0 = -2.261724623e-9
+ ua = 1.100663075e-09 lua = -5.783872961e-16
+ ub = 3.463814915e-19 lub = 2.982782283e-25
+ uc = 2.534437437e-11 luc = -6.305592823e-18 wuc = 1.938704561e-32 puc = -3.433122660e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.800738114e+04 lvsat = 1.741929099e-2
+ a0 = -2.327738550e-01 la0 = 2.058614465e-7
+ ags = 2.238513771e+00 lags = -1.772059212e-7
+ a1 = 0.0
+ a2 = 1.390223610e+00 la2 = -1.471220882e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.172705079e-02 lketa = -1.122665899e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.232093940e-01 lpclm = 2.875838254e-8
+ pdiblc1 = 4.356848163e-01 lpdiblc1 = -6.702635233e-9
+ pdiblc2 = 7.285998437e-03 lpdiblc2 = 4.754504447e-10
+ pdiblcb = -4.286388172e-01 lpdiblcb = 5.288194294e-8
+ drout = 4.877806509e-01 ldrout = 3.202728919e-10
+ pscbe1 = 7.998969111e+08 lpscbe1 = 1.848022846e-2
+ pscbe2 = 1.555222594e-08 lpscbe2 = -1.594632741e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.189402196e+00 lbeta0 = 1.912554271e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.192700175e-10 lagidl = 7.958284090e-17
+ bgidl = 1.927151494e+09 lbgidl = -1.662058126e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.636919446e-01 lkt1 = -1.338895424e-8
+ kt2 = -7.853798926e-02 lkt2 = 6.369821319e-9
+ at = 1.255074293e+05 lat = -1.332323102e-2
+ ute = -2.442725738e+00 lute = 3.934912890e-7
+ ua1 = 5.357754802e-10 lua1 = -6.115902980e-17
+ ub1 = -1.562933375e-18 lub1 = 3.462168921e-25 wub1 = 1.540743956e-39 pub1 = -3.851859889e-46
+ uc1 = -2.790687019e-10 luc1 = 4.372554830e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.89 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-3.563014349e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.429546303e-07 wvth0 = -6.015810162e-07 pvth0 = 1.180692981e-13
+ k1 = 1.177418111e+00 lk1 = -4.579641446e-08 wk1 = -1.001322624e-06 pk1 = 1.965245848e-13
+ k2 = -1.276262042e+00 lk2 = 2.235793987e-07 wk2 = 1.564647640e-06 pk2 = -3.070855691e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.079967616e+00 ldsub = -8.007548441e-07 wdsub = -2.202816395e-07 pdsub = 4.323357597e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {4.061942771e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.428541842e-07 wvoff = -6.426463607e-07 pvoff = 1.261289880e-13
+ nfactor = {1.710366912e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.852250379e-06 wnfactor = -1.761006316e-05 pnfactor = 3.456239046e-12
+ eta0 = 2.076267751e+00 leta0 = -3.274785901e-07 weta0 = -5.417325045e-07 peta0 = 1.063231300e-13
+ etab = -4.073042716e-01 letab = 7.993834622e-08 wetab = 4.837917156e-07 petab = -9.495138107e-14
+ u0 = 7.246138620e-03 lu0 = -7.022398244e-10 wu0 = -7.131486515e-09 pu0 = 1.399661201e-15
+ ua = 5.725507612e-09 lua = -1.540931844e-15 wua = -9.672579450e-15 pua = 1.898388806e-21
+ ub = -1.522754569e-20 lub = 3.975356497e-25 wub = 4.205832820e-24 pub = -8.254577784e-31
+ uc = -6.232755390e-11 luc = 1.030336826e-17 wuc = -2.129067005e-18 puc = 4.178613358e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.055251886e+06 lvsat = -3.807686012e-01 wvsat = -1.703320083e+00 pvsat = 3.343021160e-7
+ a0 = 7.405214146e+00 la0 = -1.273686083e-06 wa0 = -6.667318487e-06 pa0 = 1.308561263e-12
+ ags = 1.250000029e+00 lags = -5.611941134e-15 wags = -2.934606869e-14 pags = 5.759606125e-21
+ a1 = 0.0
+ a2 = -5.556862665e+00 la2 = 1.202395966e-06 wa2 = 4.939641162e-06 pa2 = -9.694786727e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.911848907e-01 lketa = 4.715971034e-08 wketa = -3.993273002e-08 pketa = 7.837397258e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.019473318e+00 lpclm = -6.591365094e-08 wpclm = 4.600837043e-09 ppclm = -9.029832822e-16
+ pdiblc1 = 2.193161780e+00 lpdiblc1 = -3.522694737e-07 wpdiblc1 = -4.475198705e-07 ppdiblc1 = 8.783248739e-14
+ pdiblc2 = 7.988214026e-02 lpdiblc2 = -1.372754357e-08 wpdiblc2 = -3.137794111e-08 ppdiblc2 = 6.158391612e-15
+ pdiblcb = -2.626606535e-01 lpdiblcb = 2.532112181e-08 wpdiblcb = 1.291931321e-06 ppdiblcb = -2.535609008e-13
+ drout = -2.339336619e+00 ldrout = 5.552148158e-07 wdrout = 4.419625128e-13 pdrout = -8.674177110e-20
+ pscbe1 = 7.999999956e+08 lpscbe1 = 8.667640686e-07 wpscbe1 = 4.532501221e-06 ppscbe1 = -8.895721436e-13
+ pscbe2 = -3.128838962e-08 lpscbe2 = 7.447318981e-15 wpscbe2 = 2.938289706e-14 ppscbe2 = -5.766834292e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.858738194e+01 lbeta0 = -1.831366996e-06 wbeta0 = -3.736014724e-06 pbeta0 = 7.332489297e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.943011045e-08 lagidl = 9.745495412e-15 wagidl = 4.918833966e-14 pagidl = -9.653949482e-21
+ bgidl = 9.999999969e+08 lbgidl = 6.173896790e-07 wbgidl = 3.228485107e-06 pbgidl = -6.336364746e-13
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 5.164245325e-01 lkt1 = -2.070212116e-07 wkt1 = -9.239204482e-07 pkt1 = 1.813332468e-13
+ kt2 = 2.521375380e-01 lkt2 = -5.792615022e-08 wkt2 = 5.818645121e-15 pkt2 = -1.141996497e-21
+ at = 7.784346266e+05 lat = -1.427334517e-01 wat = -5.818474433e-01 pat = 1.141962885e-7
+ ute = -2.935513576e+00 lute = 5.275237315e-07 wute = 1.378059631e-06 pute = -2.704648734e-13
+ ua1 = -2.847873369e-09 lua1 = 5.971329984e-16 wua1 = 1.375801305e-22 pua1 = -2.700216628e-29
+ ub1 = 5.029232060e-18 lub1 = -9.147621295e-25 wub1 = -7.558278787e-31 pub1 = 1.483425576e-37
+ uc1 = -1.083871809e-10 luc1 = 1.437330652e-17 wuc1 = -9.659246920e-24 puc1 = 1.895772129e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.90 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.207712395e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.065946112e-05 wvth0 = 9.447677747e-08 pvth0 = -9.447608306e-12
+ k1 = 3.837582508e-01 lk1 = 4.789700719e-06 wk1 = 4.245200426e-08 pk1 = -4.245169224e-12
+ k2 = 1.961702719e-02 lk2 = 1.946984499e-07 wk2 = 1.725648409e-09 pk2 = -1.725635725e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -2.889114370e-05 lcit = 2.921558614e-09 wcit = 2.589431491e-11 pcit = -2.589412458e-15
+ voff = {-3.615576234e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.041481379e-05 wvoff = 9.230842289e-08 pvoff = -9.230774442e-12
+ nfactor = {1.986317054e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.225829953e-07 wnfactor = -2.859112812e-09 pnfactor = 2.859091797e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.513887615e-02 lu0 = -4.630242114e-07 wu0 = -4.103869312e-09 pu0 = 4.103839148e-13
+ ua = -1.237110853e-09 lua = 4.200286056e-14 wua = 3.722791298e-16 pua = -3.722763935e-20
+ ub = 2.381952708e-18 lub = -1.142350361e-22 wub = -1.012486275e-24 pub = 1.012478833e-28
+ uc = -2.079858754e-10 luc = 1.023221334e-14 wuc = 9.069000124e-17 puc = -9.068933467e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.618781426e+05 lvsat = 2.420323636e+01 wvsat = 2.145177650e-01 pvsat = -2.145161883e-5
+ a0 = 1.928830324e+00 la0 = -4.648269077e-05 wa0 = -4.119846943e-07 pa0 = 4.119816662e-11
+ ags = -1.102248498e-01 lags = 2.235132069e-05 wags = 1.981038935e-07 pags = -1.981024375e-11
+ a1 = 0.0
+ a2 = 1.483334384e+00 la2 = -5.133306113e-05 wa2 = -4.549744248e-07 pa2 = 4.549710807e-11
+ b0 = -5.213037429e-07 lb0 = 3.916108646e-11 wb0 = 3.470919597e-13 pb0 = -3.470894086e-17
+ b1 = 2.401036046e-09 lb1 = -1.803692788e-13 wb1 = -1.598646313e-15 pb1 = 1.598634563e-19
+ keta = 9.955052647e-02 lketa = -7.618870748e-06 wketa = -6.752746203e-08 pketa = 6.752696570e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.653475026e-01 lpclm = 3.803447070e-05 wpclm = 3.371065557e-07 ppclm = -3.371040780e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 4.169528645e-03 lpdiblc2 = -2.892348586e-07 wpdiblc2 = -2.563542102e-09 ppdiblc2 = 2.563523260e-13
+ pdiblcb = -4.360120473e-01 lpdiblcb = 2.110104964e-05 wpdiblcb = 1.870225097e-07 ppdiblcb = -1.870211350e-11
+ drout = 0.56
+ pscbe1 = 8.001472062e+08 lpscbe1 = -1.472051018e+01 wpscbe1 = -1.304706071e-01 ppscbe1 = 1.304696481e-5
+ pscbe2 = 2.405702579e-08 lpscbe2 = -1.399629791e-12 wpscbe2 = -1.240517798e-14 ppscbe2 = 1.240508680e-18
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.019614025e-10 lalpha0 = 3.019591831e-14 walpha0 = 2.676320146e-16 palpha0 = -2.676300475e-20
+ alpha1 = -3.019614025e-10 lalpha1 = 3.019591831e-14 walpha1 = 2.676320146e-16 palpha1 = -2.676300475e-20
+ beta0 = 1.016295044e+02 lbeta0 = -7.162897797e-03 wbeta0 = -6.348608934e-05 pbeta0 = 6.348562272e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.294277948e-09 lagidl = -4.393988252e-13 wagidl = -3.894473140e-15 pagidl = 3.894444516e-19
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -2.271754779e+00 legidl = 2.371737347e-04 wegidl = 2.102114722e-06 pegidl = -2.102099271e-10
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.306360432e-01 lkt1 = -7.613900802e-07 wkt1 = -6.748341248e-09 pkt1 = 6.748291647e-13
+ kt2 = -7.722994633e-02 lkt2 = 1.868380900e-06 wkt2 = 1.655980584e-08 pkt2 = -1.655968412e-12
+ at = 2.853523996e+05 lat = -2.143608241e+01 wat = -1.899919672e-01 pat = 1.899905707e-5
+ ute = 6.584505920e-02 lute = -1.488239653e-05 wute = -1.319054359e-07 pute = 1.319044664e-11
+ ua1 = 2.897873375e-09 lua1 = -8.076674387e-14 wua1 = -7.158506044e-16 pua1 = 7.158453429e-20
+ ub1 = -2.777995573e-18 lub1 = 1.549084187e-22 wub1 = 1.372981995e-24 pub1 = -1.372971904e-28
+ uc1 = -9.328462329e-11 luc1 = 6.349515660e-15 wuc1 = 5.627693287e-17 puc1 = -5.627651923e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.91 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-4.140128731e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.213945940e-06 wvth0 = -6.298451831e-07 pvth0 = 5.038298529e-12
+ k1 = 7.403975898e-01 lk1 = -2.342823932e-06 wk1 = -2.830133617e-07 pk1 = 2.263898879e-12
+ k2 = 3.411420156e-02 lk2 = -9.523438199e-08 wk2 = -1.150432273e-08 pk2 = 9.202612613e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.886470271e-04 lcit = -1.429044911e-09 wcit = -1.726287660e-10 pcit = 1.380903246e-15
+ voff = {4.139255487e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.094279669e-06 wvoff = -6.153894859e-07 pvoff = 4.922663576e-12
+ nfactor = {1.962297643e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.577875541e-07 wnfactor = 1.906075208e-08 pnfactor = -1.524720070e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = -1.933773489e-02 lu0 = 2.264826692e-07 wu0 = 2.735912874e-08 pu0 = -2.188529210e-13
+ ua = 1.890406566e-09 lua = -2.054518908e-14 wua = -2.481860865e-15 pua = 1.985306275e-20
+ ub = -6.123945712e-18 lub = 5.587668043e-23 wub = 6.749908501e-24 pub = -5.399430682e-29
+ uc = 5.539009345e-10 luc = -5.004962875e-15 wuc = -6.046000083e-16 puc = 4.836355685e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.640285860e+06 lvsat = -1.183871910e+01 wvsat = -1.430118433e+00 pvsat = 1.143989633e-5
+ a0 = -1.532253590e+00 la0 = 2.273644362e-05 wa0 = 2.746564629e-06 pa0 = -2.197049830e-11
+ ags = 1.554046199e+00 lags = -1.093287704e-05 wags = -1.320692623e-06 pags = 1.056457028e-11
+ a1 = 0.0
+ a2 = -2.338906308e+00 la2 = 2.510894336e-05 wa2 = 3.033162832e-06 pa2 = -2.426307328e-11
+ b0 = 2.394616230e-06 lb0 = -1.915516979e-11 wb0 = -2.313946398e-12 pb0 = 1.850987043e-17
+ b1 = -1.102919356e-08 lb1 = 8.822544200e-14 wb1 = 1.065764208e-14 pb1 = -8.525330331e-20
+ keta = -4.677477636e-01 lketa = 3.726678088e-06 wketa = 4.501830802e-07 pketa = -3.601133757e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.466685079e+00 lpclm = -1.860409938e-05 wpclm = -2.247377038e-06 ppclm = 1.797736448e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -1.736679165e-02 lpdiblc2 = 1.414757181e-07 wpdiblc2 = 1.709028068e-08 ppdiblc2 = -1.367096841e-13
+ pdiblcb = 1.135164282e+00 lpdiblcb = -1.032132214e-05 wpdiblcb = -1.246816731e-06 ppdiblcb = 9.973617438e-12
+ drout = 0.56
+ pscbe1 = 7.990511225e+08 lpscbe1 = 7.200358759e+00 wpscbe1 = 8.698040474e-01 ppscbe1 = -6.957793073e-6
+ pscbe2 = -8.015888936e-08 lpscbe2 = 6.846119127e-13 wpscbe2 = 8.270118650e-14 ppscbe2 = -6.615487066e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.946415475e-09 lalpha0 = -1.476996669e-14 walpha0 = -1.784213431e-15 palpha0 = 1.427239605e-20
+ alpha1 = 1.946415475e-09 lalpha1 = -1.476996669e-14 walpha1 = -1.784213431e-15 palpha1 = 1.427239605e-20
+ beta0 = -4.317172088e+02 lbeta0 = 3.503644458e-03 wbeta0 = 4.232405956e-04 pbeta0 = -3.385613683e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.642319560e-08 lagidl = 2.149265985e-13 wagidl = 2.596315427e-14 pagidl = -2.076861512e-19
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.538811354e+01 legidl = -1.160106516e-04 wegidl = -1.401409815e-05 pegidl = 1.121024848e-10
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.873288662e-01 lkt1 = 3.724247100e-07 wkt1 = 4.498894165e-08 pkt1 = -3.598784663e-13
+ kt2 = 6.188900252e-02 lkt2 = -9.138958242e-07 wkt2 = -1.103987056e-07 pkt2 = 8.831085017e-13
+ at = -1.310770346e+06 lat = 1.048519935e+01 wat = 1.266613114e+00 pat = -1.013197395e-5
+ ute = -1.042292667e+00 lute = 7.279543504e-06 wute = 8.793695724e-07 pute = -7.034310243e-12
+ ua1 = -3.115988417e-09 lua1 = 3.950607178e-14 wua1 = 4.772337363e-15 pua1 = -3.817519123e-20
+ ub1 = 8.756427829e-18 lub1 = -7.577157152e-23 wub1 = -9.153213303e-24 pub1 = 7.321897881e-29
+ uc1 = 3.794979577e-10 luc1 = -3.105788465e-15 wuc1 = -3.751795525e-16 puc1 = 3.001160663e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.92 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.069866256e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.239906809e-8
+ k1 = 4.556237202e-01 lk1 = -6.484228401e-8
+ k2 = 2.007683582e-02 lk2 = 1.705422642e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.164179846e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.199470589e-8
+ nfactor = {2.378038919e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.167837078e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.443397737e-03 lu0 = 4.254027232e-9
+ ua = -7.572954228e-10 lua = 6.344807637e-16 wua = 1.654361225e-30
+ ub = 8.922232633e-19 lub = -2.475144842e-25
+ uc = -7.084368051e-11 luc = -7.465141979e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.671623623e+05 lvsat = -8.547403617e-1
+ a0 = 1.370094967e+00 la0 = -4.802116133e-7
+ ags = 1.321801322e-01 lags = 4.410064215e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.426888399e-04 lketa = -8.219334060e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.401119263e-01 lpclm = -7.931506930e-07 ppclm = 1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.387319811e-03 lpdiblc2 = 1.365168829e-08 ppdiblc2 = -1.387778781e-29
+ pdiblcb = -2.488330300e-01 lpdiblcb = 7.496391204e-07 ppdiblcb = -1.776356839e-27
+ drout = 0.56
+ pscbe1 = 1.224636900e+09 lpscbe1 = -3.397173053e+3
+ pscbe2 = -1.698011262e-08 lpscbe2 = 1.792281353e-13 ppscbe2 = 2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.446751046e+00 lbeta0 = 2.265262463e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.904539975e-10 lagidl = -1.962669803e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.670754974e+00 legidl = -6.281865390e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.063193317e-01 lkt1 = -2.755920237e-7
+ kt2 = -4.841666844e-02 lkt2 = -3.153153126e-8
+ at = -9.065933829e+04 lat = 7.252080717e-1
+ ute = -1.645263111e-01 lute = 2.580578176e-7
+ ua1 = 5.778773827e-10 lua1 = 9.957860376e-15
+ ub1 = 8.146409535e-19 lub1 = -1.224311373e-23
+ uc1 = -1.163111597e-11 luc1 = 2.295664482e-17 wuc1 = -2.584939414e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.93 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063199473e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.736836213e-9
+ k1 = 4.427665361e-01 lk1 = -1.342299740e-8
+ k2 = 2.238297990e-02 lk2 = 7.831345119e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.585912374e-01 ldsub = -1.194145485e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.482687602e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.538498620e-8
+ nfactor = {9.059919706e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.719268760e-6
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394757071e-01 letab = 2.778517638e-7
+ u0 = 8.601632881e-03 lu0 = 3.621202956e-9
+ ua = -7.352853466e-10 lua = 5.464566366e-16
+ ub = 8.528601283e-19 lub = -9.009087610e-26
+ uc = -7.556913799e-11 luc = 1.143321474e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.264314745e+00 la0 = -5.716847236e-8
+ ags = 1.560797535e-01 lags = 3.454255025e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.464757958e-03 lketa = -3.744375028e-08 wketa = 6.938893904e-24 pketa = -2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.488073345e-01 lpclm = 2.361946495e-06 wpclm = -1.110223025e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 3.621872386e-03 lpdiblc2 = -6.381398745e-9
+ pdiblcb = -9.776424111e-02 lpdiblcb = 1.454750005e-7
+ drout = 0.56
+ pscbe1 = -4.171210305e+07 lpscbe1 = 1.667292191e+3
+ pscbe2 = 4.631193739e-08 lpscbe2 = -7.389354511e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.144527102e+01 lbeta0 = -9.335576356e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.690680066e-10 lagidl = -2.774355581e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815376811e-01 lkt1 = 2.522608815e-8
+ kt2 = -6.023855242e-02 lkt2 = 1.574731557e-8
+ at = 1.021557796e+05 lat = -4.591068088e-2
+ ute = -1.323451088e-01 lute = 1.293566616e-7
+ ua1 = 3.320607059e-09 lua1 = -1.011042424e-15
+ ub1 = -2.835183653e-18 lub1 = 2.353502076e-24
+ uc1 = 1.789645493e-11 luc1 = -9.513193603e-17 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.94 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.080253346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.983204748e-8
+ k1 = 3.559763493e-01 lk1 = 1.600935854e-7
+ k2 = 5.664373486e-02 lk2 = -6.066498314e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.538016126e-01 ldsub = 1.029822606e-06 pdsub = 8.881784197e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.107617634e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.985602103e-10
+ nfactor = {2.269123695e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.992787282e-9
+ eta0 = -2.188386675e-01 leta0 = 4.385161211e-07 weta0 = -1.457167720e-22 peta0 = -7.112366252e-29
+ etab = 8.242798594e-01 letab = -1.648951009e-06 wetab = 4.423544864e-22 petab = -4.024558464e-28
+ u0 = 1.231769894e-02 lu0 = -3.808197859e-9
+ ua = -2.809317911e-10 lua = -3.619165246e-16
+ ub = 9.337272840e-19 lub = -2.517657501e-25
+ uc = -7.496753916e-11 luc = 1.023045924e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.949154737e+04 lvsat = -1.210264538e-2
+ a0 = 1.349266482e+00 la0 = -2.270095072e-7
+ ags = 1.615750419e-01 lags = 3.344389646e-7
+ a1 = 0.0
+ a2 = 6.001569927e-01 la2 = 3.995391301e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.083405179e-02 lketa = -2.858845418e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.592302506e-01 lpclm = 3.466122321e-7
+ pdiblc1 = 7.407420150e-01 lpdiblc1 = -7.012262346e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.203234000e-01 ldrout = 8.790300377e-7
+ pscbe1 = 7.981743154e+08 lpscbe1 = -1.186332945e+1
+ pscbe2 = 9.526279703e-09 lpscbe2 = -3.492672025e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.883960260e+00 lbeta0 = 1.782957602e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.471808281e-10 lagidl = 7.546826683e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.587827164e-01 lkt1 = -2.026711633e-8
+ kt2 = -5.616202393e-02 lkt2 = 7.597254838e-9
+ at = 9.660944576e+04 lat = -3.482208970e-2
+ ute = 9.121531202e-01 lute = -1.958872090e-06 pute = -2.220446049e-28
+ ua1 = 6.057818692e-09 lua1 = -6.483453838e-15 pua1 = -1.323488980e-35
+ ub1 = -4.209009179e-18 lub1 = 5.100143366e-24 pub1 = 6.162975822e-45
+ uc1 = -1.262217768e-10 luc1 = 1.929986004e-16 wuc1 = -1.033975766e-31 puc1 = 1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.95 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.090058366e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.962986083e-08 wvth0 = 2.540412968e-08 pvth0 = -2.538545764e-14
+ k1 = 4.467888797e-01 lk1 = 6.934780215e-08 wk1 = 6.720919733e-08 pk1 = -6.715979857e-14
+ k2 = 1.227178436e-03 lk2 = -5.289157886e-09 wk2 = -6.179796102e-09 pk2 = 6.175253952e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.922799802e+00 ldsub = -1.145179006e-06 wdsub = -6.112380655e-07 pdsub = 6.107888055e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {4.655183889e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.567259166e-07 wvoff = -2.299290755e-07 pvoff = 2.297600777e-13
+ nfactor = {-5.249657284e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.507261888e-06 wnfactor = 6.821426369e-06 pnfactor = -6.816412621e-12
+ eta0 = -4.628912179e-01 leta0 = 6.823892929e-07 weta0 = 3.993652678e-07 peta0 = -3.990717344e-13
+ etab = -1.650251575e+00 letab = 8.237616446e-07 wetab = 3.108292652e-10 petab = -3.106008057e-16
+ u0 = -1.347251501e-02 lu0 = 2.196306029e-08 wu0 = 2.113707965e-08 pu0 = -2.112154390e-14
+ ua = -6.102674040e-09 lua = 5.455546744e-15 wua = 5.332260492e-15 pua = -5.328341281e-21
+ ub = 4.062452390e-18 lub = -3.378191243e-24 wub = -3.486976601e-24 pub = 3.484413674e-30
+ uc = -1.156356345e-10 luc = 5.086866353e-17 wuc = 1.541949103e-17 puc = -1.540815770e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.320865357e+05 lvsat = -6.842032764e-01 wvsat = -6.681545105e-01 pvsat = 6.676634169e-7
+ a0 = 1.868314391e+00 la0 = -7.456759162e-07 wa0 = -3.297255827e-07 pa0 = 3.294832344e-13
+ ags = -2.563720029e-01 lags = 7.520788183e-07 wags = 6.314557766e-16 pags = -6.309930356e-22
+ a1 = 0.0
+ a2 = 5.827741276e-01 la2 = 4.169092188e-07 wa2 = 4.127133425e-07 pa2 = -4.124099982e-13
+ b0 = 9.702731453e-16 lb0 = -9.695599945e-22 wb0 = -9.375865836e-22 pb0 = 9.368974574e-28
+ b1 = 4.033869646e-19 lb1 = -4.030904751e-25 wb1 = -3.897976645e-25 pb1 = 3.895111632e-31
+ keta = 5.306598703e-03 lketa = -1.898763253e-08 wketa = 4.818116172e-09 pketa = -4.814574856e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.930301530e+00 lpclm = -1.123377810e-06 wpclm = -3.354036300e-07 ppclm = 3.351571083e-13
+ pdiblc1 = 1.174558853e-01 lpdiblc1 = -7.839822018e-08 wpdiblc1 = -4.879617772e-08 ppdiblc1 = 4.876031252e-14
+ pdiblc2 = 1.474177464e-03 lpdiblc2 = -1.043409994e-09 wpdiblc2 = -6.328242120e-10 ppdiblc2 = 6.323590862e-16
+ pdiblcb = -2.067049663e-01 lpdiblcb = 1.815714132e-07 wpdiblcb = 1.703049107e-07 ppdiblcb = -1.701797366e-13
+ drout = 5.813977084e-01 ldrout = 4.182946189e-07 wdrout = 4.045004176e-07 pdrout = -4.042031098e-13
+ pscbe1 = 2.050399128e+08 lpscbe1 = 5.808351193e+02 wpscbe1 = 5.484639480e+02 ppscbe1 = -5.480608270e-4
+ pscbe2 = 6.807869009e-08 lpscbe2 = -5.885864157e-14 wpscbe2 = -5.706372530e-14 ppscbe2 = 5.702178346e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.321044596e+00 lbeta0 = 1.346194523e-06 wbeta0 = 2.564908231e-07 pbeta0 = -2.563023023e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.307246020e-09 lagidl = 1.813968712e-15 wagidl = 2.058559823e-15 pagidl = -2.057046781e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.736648681e-01 lkt1 = -1.053224030e-07 wkt1 = -4.491548589e-08 pkt1 = 4.488247301e-14
+ kt2 = -8.748539788e-02 lkt2 = 3.889760611e-08 wkt2 = 2.227871000e-08 pkt2 = -2.226233515e-14
+ at = 1.269138733e+05 lat = -6.510424351e-02 wat = -3.722291157e-02 pat = 3.719555273e-8
+ ute = -1.930873461e+00 lute = 8.820648669e-07 wute = 3.319551114e-08 pute = -3.317111244e-14
+ ua1 = -4.195647473e-09 lua1 = 3.762476029e-15 wua1 = 7.467127104e-16 pua1 = -7.461638766e-22
+ ub1 = 5.571987544e-18 lub1 = -4.673664324e-24 wub1 = -1.303087838e-24 pub1 = 1.302130068e-30
+ uc1 = 4.385574696e-10 luc1 = -3.713655331e-16 wuc1 = -1.060772972e-16 puc1 = 1.059993304e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.96 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.175937290e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.250620212e-08 wvth0 = 1.532371786e-07 pvth0 = -8.920802483e-14
+ k1 = 1.093389577e+00 lk1 = -2.534772949e-07 wk1 = -5.774850110e-07 pk1 = 2.547134553e-13
+ k2 = -2.802008634e-01 lk2 = 1.352180134e-07 wk2 = 2.585888821e-07 pk2 = -1.260144802e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.877967906e+00 ldsub = 7.524112834e-07 wdsub = 1.537040934e-06 pdsub = -4.617717091e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-8.225677897e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.771950948e-07 wvoff = 5.744974259e-07 pvoff = -1.718619196e-13
+ nfactor = {1.753731822e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.869477435e-06 wnfactor = -1.421958829e-05 pnfactor = 3.688629565e-12
+ eta0 = 1.316576242e+00 leta0 = -2.060365284e-07 weta0 = -7.987305414e-07 peta0 = 1.990955698e-13
+ etab = -1.322736607e-03 letab = 5.091882339e-10 wetab = 7.808354845e-11 petab = -1.943990154e-16
+ u0 = 4.976590408e-02 lu0 = -9.609669019e-09 wu0 = -3.841768815e-08 pu0 = 8.612067246e-15
+ ua = 9.917435451e-09 lua = -2.542733221e-15 wua = -9.762500269e-15 pua = 2.207944451e-21
+ ub = -6.432634963e-18 lub = 1.861638544e-24 wub = 6.485342485e-24 pub = -1.494416215e-30
+ uc = -3.896393326e-11 luc = 1.258916661e-17 wuc = -1.976524315e-17 puc = 2.158348607e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.245401567e+06 lvsat = 3.030873212e-01 wvsat = 1.223228867e+00 pvsat = -2.766381049e-7
+ a0 = 4.040946006e-01 la0 = -1.464222245e-08 wa0 = 4.207541152e-07 pa0 = -4.520501195e-14
+ ags = 7.317898639e-01 lags = 2.587241839e-07 wags = 2.332931116e-07 pags = -1.164750857e-13
+ a1 = 0.0
+ a2 = 1.989880832e+00 la2 = -2.856099102e-07 wa2 = -7.829640928e-07 pa2 = 1.845498966e-13
+ b0 = -1.940546291e-15 lb0 = 4.837102711e-22 wb0 = 1.875173167e-21 pb0 = -4.674150395e-28
+ b1 = -8.067739291e-19 lb1 = 2.011005034e-25 wb1 = 7.795953290e-25 pb1 = -1.943258297e-31
+ keta = -1.408755808e-02 lketa = -9.304808842e-09 wketa = -2.707943301e-08 pketa = 1.111075503e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.290542050e+00 lpclm = 4.846766597e-07 wpclm = 6.855474741e-07 ppclm = -1.745680447e-13
+ pdiblc1 = -5.326323903e-01 lpdiblc1 = 2.461681027e-07 wpdiblc1 = 1.420548808e-07 ppdiblc1 = -4.652494118e-14
+ pdiblc2 = -1.721043617e-02 lpdiblc2 = 8.285163633e-09 wpdiblc2 = 7.850521310e-09 ppdiblc2 = -3.603078416e-15
+ pdiblcb = -2.608375325e-01 lpdiblcb = 2.085979089e-07 wpdiblcb = 4.229426830e-07 ppdiblcb = -2.963129340e-13
+ drout = 2.784244617e+00 ldrout = -6.815097430e-07 wdrout = -1.231866408e-06 pdrout = 4.127775735e-13
+ pscbe1 = 1.935223156e+09 lpscbe1 = -2.829848175e+02 wpscbe1 = -1.096951866e+03 ppscbe1 = 2.734376992e-4
+ pscbe2 = -1.120315279e-07 lpscbe2 = 3.106408640e-14 wpscbe2 = 1.174382471e-13 ppscbe2 = -3.010094380e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.561703869e+00 lbeta0 = 2.275117714e-07 wbeta0 = -1.414000253e-08 pbeta0 = -1.211858032e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.453239534e-09 lagidl = -5.627751077e-16 wagidl = -3.061635815e-15 pagidl = 4.992876940e-22
+ bgidl = 5.139579501e+08 lbgidl = 2.426637841e+02 wbgidl = 2.188113332e+02 pbgidl = -1.092448403e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.118922597e-01 lkt1 = 6.354269570e-08 wkt1 = 1.480570615e-07 pkt1 = -5.146196586e-14
+ kt2 = 3.558679744e-02 lkt2 = -2.254803349e-08 wkt2 = -4.637617321e-08 pkt2 = 1.201464512e-14
+ at = -1.248673637e+05 lat = 6.060131579e-02 wat = 1.189536670e-01 pat = -4.077794677e-8
+ ute = 8.599772217e-01 lute = -5.113091994e-07 wute = -3.816106357e-07 pute = 1.739270785e-13
+ ua1 = 6.432394267e-09 lua1 = -1.543733230e-15 wua1 = -1.542720933e-15 pua1 = 3.968702112e-22
+ ub1 = -7.342107914e-18 lub1 = 1.773891545e-24 wub1 = 2.556424953e-24 pub1 = -6.247895851e-31
+ uc1 = -4.426110368e-10 luc1 = 6.857106122e-17 wuc1 = 1.506203596e-16 puc1 = -2.216082522e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.97 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.006168271e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.387844688e-08 wvth0 = 5.638090250e-08 pvth0 = -6.506514516e-14
+ k1 = 2.582520869e+00 lk1 = -6.246656064e-07 wk1 = -2.986207367e-06 pk1 = 8.551236334e-13
+ k2 = -1.191749899e+00 lk2 = 3.624352838e-07 wk2 = 1.513914113e-06 pk2 = -4.389231238e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.808340898e+01 ldsub = 4.791860552e-06 wdsub = 1.780071519e-05 pdsub = -4.515736473e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {4.974656646e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.518430442e-07 wvoff = -4.784590195e-07 pvoff = 9.060326879e-14
+ nfactor = {3.025313879e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.039086451e-06 wnfactor = -2.660727576e-05 pnfactor = 6.776446482e-12
+ eta0 = -4.639882971e+00 leta0 = 1.278700277e-06 weta0 = 5.160695607e-06 peta0 = -1.286380789e-12
+ etab = -7.737488982e-01 letab = 1.930479954e-07 wetab = 7.476768058e-07 petab = -1.865445945e-13
+ u0 = 7.587355088e-02 lu0 = -1.611739160e-08 wu0 = -5.758134939e-08 pu0 = 1.338889727e-14
+ ua = 2.139979803e-08 lua = -5.404884329e-15 wua = -1.961529769e-14 pua = 4.663902001e-21
+ ub = -1.594397075e-17 lub = 4.232481658e-24 wub = 1.574156285e-23 pub = -3.801667985e-30
+ uc = 3.476162990e-10 luc = -8.377175499e-17 wuc = -3.114152280e-16 puc = 7.485648209e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.605410077e+06 lvsat = 3.928248424e-01 wvsat = 1.568727771e+00 pvsat = -3.627588892e-7
+ a0 = 5.061943530e+00 la0 = -1.175680936e-06 wa0 = -5.116348946e-06 pa0 = 1.335000983e-12
+ ags = 3.100750734e+00 lags = -3.317748473e-07 wags = -8.331899237e-07 pags = 1.493618081e-13
+ a1 = 0.0
+ a2 = 3.694349257e+00 la2 = -7.104742321e-07 wa2 = -2.226504262e-06 pa2 = 5.443739369e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.413342252e+00 lketa = -3.651131005e-07 wketa = -1.354397589e-06 pketa = 3.419647151e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.168805833e+00 lpclm = 4.543320817e-07 wpclm = 1.635014618e-06 ppclm = -4.112369724e-13
+ pdiblc1 = -5.941634316e+00 lpdiblc1 = 1.594442968e-06 wpdiblc1 = 6.162480006e-06 ppdiblc1 = -1.547206210e-12
+ pdiblc2 = -1.408564542e-01 lpdiblc2 = 3.910578831e-08 wpdiblc2 = 1.431518297e-07 ppdiblc2 = -3.732895905e-14
+ pdiblcb = -4.587364896e+00 lpdiblcb = 1.287049752e-06 wpdiblcb = 4.018626914e-06 ppdiblcb = -1.192591164e-12
+ drout = 1.340703730e+01 ldrout = -3.329400162e-06 wdrout = -1.248403273e-05 pdrout = 3.217548812e-12
+ pscbe1 = 7.998083225e+08 lpscbe1 = 3.436096044e-02 wpscbe1 = 8.560428009e-02 ppscbe1 = -1.534574189e-8
+ pscbe2 = 4.825581032e-08 lpscbe2 = -8.889936954e-15 wpscbe2 = -3.160186603e-14 ppscbe2 = 7.049540005e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -1.563904373e+01 lbeta0 = 6.259911123e-06 wbeta0 = 2.302571324e-05 pbeta0 = -5.864214823e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.813022266e-09 lagidl = -6.524563505e-16 wagidl = -3.896452421e-15 pagidl = 7.073782551e-22
+ bgidl = 2.735865702e+09 lbgidl = -3.111800517e+02 wbgidl = -7.814702435e+02 pbgidl = 1.400903469e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.886265556e-01 lkt1 = -6.688913004e-08 wkt1 = -2.657989862e-07 pkt1 = 5.169786187e-14
+ kt2 = -1.596197014e+00 lkt2 = 3.841985582e-07 wkt2 = 1.466532127e-06 pkt2 = -3.651004424e-13
+ at = 8.354122558e+03 lat = 2.739386202e-02 wat = 1.132066461e-01 pat = -3.934541561e-8
+ ute = 2.001439250e+00 lute = -7.958357319e-07 wute = -4.294449958e-06 pute = 1.149260972e-12
+ ua1 = 1.592910468e-08 lua1 = -3.910930751e-15 wua1 = -1.487475872e-14 pua1 = 3.720080611e-21
+ ub1 = -2.560732494e-17 lub1 = 6.326770866e-24 wub1 = 2.323438410e-23 pub1 = -5.779081072e-30
+ uc1 = -1.315842322e-10 luc1 = -8.957035249e-18 wuc1 = -1.425160129e-16 puc1 = 5.090781267e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.98 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {6.892783141e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.858978899e-07 wvth0 = -1.611937275e-06 pvth0 = 2.561970853e-13
+ k1 = -1.089284020e+01 lk1 = 1.960838049e-06 wk1 = 1.066231283e-05 pk1 = -1.742510377e-12
+ k2 = 6.257877035e+00 lk2 = -1.065295402e-06 wk2 = -5.715681360e-06 pk2 = 9.383696172e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.511081367e+01 ldsub = -9.119183398e-06 wdsub = -4.856568855e-05 pdsub = 8.081430909e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {2.236942682e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.125108311e-07 wvoff = -4.662944121e-07 pvoff = 9.680784174e-14
+ nfactor = {-5.868245665e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.748329839e-06 wnfactor = 5.562297961e-05 pnfactor = -8.719852826e-12
+ eta0 = 1.571828722e+01 leta0 = -2.595634708e-06 weta0 = -1.372417962e-05 peta0 = 2.298069604e-12
+ etab = 1.572254645e+00 letab = -2.490833255e-07 wetab = -1.429079820e-06 petab = 2.229862086e-13
+ u0 = -8.224266013e-02 lu0 = 1.338684733e-08 wu0 = 7.934261358e-08 pu0 = -1.221479279e-14
+ ua = -3.761421063e-08 lua = 5.664945853e-15 wua = 3.220711037e-14 pua = -5.064737284e-21
+ ub = 3.698697261e-17 lub = -5.754636619e-24 wub = -3.154983721e-23 pub = 5.119460111e-30
+ uc = -7.810350828e-10 luc = 1.297987927e-16 wuc = 6.923666427e-16 puc = -1.150520013e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.381868750e+06 lvsat = -5.487511992e-01 wvsat = -2.985245878e+00 pvsat = 4.966257162e-7
+ a0 = -8.374408238e+00 la0 = 1.349912853e-06 wa0 = 8.580719978e-06 pa0 = -1.226653872e-12
+ ags = 1.249999377e+00 lags = 1.036146884e-13 wags = 6.001708215e-13 pags = -9.978740323e-20
+ a1 = 0.0
+ a2 = -1.107941345e+01 la2 = 2.121722845e-06 wa2 = 1.027614826e-05 pa2 = -1.857835268e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.036454107e+00 lketa = 6.698668956e-07 wketa = 3.579165857e-06 pketa = -5.938920283e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.481045060e+00 lpclm = -8.077158321e-07 wpclm = -4.306669476e-06 ppclm = 7.159093660e-13
+ pdiblc1 = 1.890788987e+01 lpdiblc1 = -3.131445200e-06 wpdiblc1 = -1.659916220e-05 ppdiblc1 = 2.773383342e-12
+ pdiblc2 = 5.207372550e-01 lpdiblc2 = -8.703343367e-08 wpdiblc2 = -4.573815288e-07 ppdiblc2 = 7.699475289e-14
+ pdiblcb = 1.756069672e+01 lpdiblcb = -2.937786479e-06 wpdiblcb = -1.593099279e-05 ppdiblcb = 2.609725531e-12
+ drout = -3.933551919e+01 ldrout = 6.706385099e-06 wdrout = 3.574985562e-05 pdrout = -5.943949745e-12
+ pscbe1 = 7.999999961e+08 lpscbe1 = 6.330432892e-07 wpscbe1 = 3.991966248e-06 ppscbe1 = -6.637248993e-13
+ pscbe2 = -8.379582697e-08 lpscbe2 = 1.618413004e-14 wpscbe2 = 8.012146386e-14 ppscbe2 = -1.420931966e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.419783570e+01 lbeta0 = -1.274093617e-05 wbeta0 = -6.713618352e-05 pbeta0 = 1.127529654e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.153500980e-09 lagidl = -1.923589331e-16 wagidl = 3.087889300e-16 pagidl = -5.088157469e-23
+ bgidl = 9.999968377e+08 lbgidl = 5.257670002e-04 wbgidl = 3.055916809e-03 pbgidl = -5.080920048e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 3.615447546e-01 lkt1 = -1.812117104e-07 wkt1 = -7.742582602e-07 pkt1 = 1.563932160e-13
+ kt2 = 4.111988207e+00 lkt2 = -6.996842218e-07 wkt2 = -3.729820014e-06 pkt2 = 6.201385245e-13
+ at = 1.502341063e+06 lat = -2.632256790e-01 wat = -1.281366920e+00 pat = 2.306293736e-7
+ ute = -1.727522377e+01 lute = 2.912028102e-06 wute = 1.523469367e-05 pute = -2.574640060e-12
+ ua1 = -4.263721532e-08 lua1 = 7.212707935e-15 wua1 = 3.844891874e-14 pua1 = -6.392709475e-21
+ ub1 = 6.598347822e-17 lub1 = -1.104931985e-23 wub1 = -5.890082027e-23 pub1 = 9.793144884e-30
+ uc1 = -1.066137913e-09 luc1 = 1.736137323e-16 wuc1 = 9.254860159e-16 puc1 = -1.538759324e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.99 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.100 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.124648838e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.706194604e-7
+ k1 = 4.210818616e-01 lk1 = 2.114671972e-7
+ k2 = 2.113420949e-02 lk2 = 8.596014224e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = 1.016439537e-26 pcit = -1.355252716e-31
+ voff = {-2.804004741e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.598181832e-7
+ nfactor = {1.983803335e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.424216791e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.153077275e-02 lu0 = -2.044270362e-8
+ ua = -9.098047201e-10 lua = 1.854443048e-15
+ ub = 1.491779338e-18 lub = -5.043522411e-24
+ uc = -1.282516351e-10 luc = 4.517563002e-16 wuc = -8.271806126e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.672490943e+04 lvsat = 1.068582539e+0
+ a0 = 1.566615238e+00 la0 = -2.052229338e-6
+ ags = 6.394720045e-02 lags = 9.868197240e-7
+ a1 = 0.0
+ a2 = 1.083322921e+00 la2 = -2.266375124e-6
+ b0 = -2.161420565e-07 lb0 = 1.728977587e-12
+ b1 = 9.955134135e-10 lb1 = -7.963375606e-15
+ keta = 4.018068624e-02 lketa = -3.363761825e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.896493835e-02 lpclm = 1.679237053e-06 ppclm = -2.664535259e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.915673984e-03 lpdiblc2 = -1.276983438e-8
+ pdiblcb = -2.715826998e-01 lpdiblcb = 9.316197581e-7
+ drout = 0.56
+ pscbe1 = 8.000324970e+08 lpscbe1 = -6.499163960e-1
+ pscbe2 = 1.315044923e-08 lpscbe2 = -6.179421357e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.666054167e-11 lalpha0 = 1.333161838e-15
+ alpha1 = -6.666054167e-11 lalpha1 = 1.333161838e-15
+ beta0 = 4.581282086e+01 lbeta0 = -3.162447948e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.870274718e-09 lagidl = -1.939963340e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.235849912e-01 legidl = 1.047131499e-05 pegidl = 7.105427358e-27
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365691544e-01 lkt1 = -3.361567574e-8
+ kt2 = -6.267063968e-02 lkt2 = 8.248976200e-8
+ at = 1.183123185e+05 lat = -9.464115887e-1
+ ute = -5.012560544e-02 lute = -6.570637432e-7
+ ua1 = 2.268500750e-09 lua1 = -3.565883958e-15
+ ub1 = -1.570875991e-18 lub1 = 6.839268476e-24
+ uc1 = -4.380619758e-11 luc1 = 2.803336491e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.101 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.069866256e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.239906809e-8
+ k1 = 4.556237202e-01 lk1 = -6.484228401e-8
+ k2 = 2.007683582e-02 lk2 = 1.705422642e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.164179846e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.199470589e-8
+ nfactor = {2.378038919e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.167837078e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.443397737e-03 lu0 = 4.254027232e-9
+ ua = -7.572954228e-10 lua = 6.344807637e-16
+ ub = 8.922232633e-19 lub = -2.475144842e-25
+ uc = -7.084368051e-11 luc = -7.465141979e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.671623623e+05 lvsat = -8.547403617e-1
+ a0 = 1.370094967e+00 la0 = -4.802116133e-7
+ ags = 1.321801322e-01 lags = 4.410064215e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.426888399e-04 lketa = -8.219334060e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.401119263e-01 lpclm = -7.931506930e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.387319811e-03 lpdiblc2 = 1.365168829e-08 ppdiblc2 = -2.775557562e-29
+ pdiblcb = -2.488330300e-01 lpdiblcb = 7.496391204e-7
+ drout = 0.56
+ pscbe1 = 1.224636900e+09 lpscbe1 = -3.397173053e+3
+ pscbe2 = -1.698011262e-08 lpscbe2 = 1.792281353e-13 ppscbe2 = 2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.446751046e+00 lbeta0 = 2.265262463e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.904539975e-10 lagidl = -1.962669803e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.670754974e+00 legidl = -6.281865390e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.063193317e-01 lkt1 = -2.755920237e-7
+ kt2 = -4.841666844e-02 lkt2 = -3.153153126e-8
+ at = -9.065933829e+04 lat = 7.252080717e-1
+ ute = -1.645263111e-01 lute = 2.580578176e-7
+ ua1 = 5.778773827e-10 lua1 = 9.957860376e-15
+ ub1 = 8.146409535e-19 lub1 = -1.224311373e-23 pub1 = -2.465190329e-44
+ uc1 = -1.163111597e-11 luc1 = 2.295664482e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.102 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063199473e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.736836213e-9
+ k1 = 4.427665361e-01 lk1 = -1.342299740e-8
+ k2 = 2.238297990e-02 lk2 = 7.831345119e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.585912374e-01 ldsub = -1.194145485e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.482687602e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.538498620e-8
+ nfactor = {9.059919706e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.719268760e-6
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394757071e-01 letab = 2.778517638e-7
+ u0 = 8.601632882e-03 lu0 = 3.621202956e-9
+ ua = -7.352853466e-10 lua = 5.464566366e-16
+ ub = 8.528601283e-19 lub = -9.009087610e-26
+ uc = -7.556913799e-11 luc = 1.143321474e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.264314745e+00 la0 = -5.716847236e-8
+ ags = 1.560797535e-01 lags = 3.454255025e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.464757958e-03 lketa = -3.744375028e-08 pketa = -5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.488073345e-01 lpclm = 2.361946495e-06 wpclm = -8.881784197e-22 ppclm = -4.440892099e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.621872386e-03 lpdiblc2 = -6.381398745e-9
+ pdiblcb = -9.776424111e-02 lpdiblcb = 1.454750005e-7
+ drout = 0.56
+ pscbe1 = -4.171210305e+07 lpscbe1 = 1.667292191e+3
+ pscbe2 = 4.631193739e-08 lpscbe2 = -7.389354511e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.144527102e+01 lbeta0 = -9.335576356e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.690680066e-10 lagidl = -2.774355581e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815376811e-01 lkt1 = 2.522608815e-8
+ kt2 = -6.023855242e-02 lkt2 = 1.574731557e-8
+ at = 1.021557796e+05 lat = -4.591068088e-2
+ ute = -1.323451088e-01 lute = 1.293566616e-7
+ ua1 = 3.320607059e-09 lua1 = -1.011042424e-15 wua1 = 2.646977960e-29
+ ub1 = -2.835183653e-18 lub1 = 2.353502076e-24
+ uc1 = 1.789645493e-11 luc1 = -9.513193603e-17 wuc1 = -5.169878828e-32 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.103 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.080253346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.983204748e-8
+ k1 = 3.559763493e-01 lk1 = 1.600935854e-7
+ k2 = 5.664373486e-02 lk2 = -6.066498314e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.538016126e-01 ldsub = 1.029822606e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.107617634e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.985602103e-10
+ nfactor = {2.269123695e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.992787282e-9
+ eta0 = -2.188386675e-01 leta0 = 4.385161211e-07 weta0 = -7.563394355e-22 peta0 = 1.401656569e-27
+ etab = 8.242798594e-01 letab = -1.648951009e-06 wetab = 1.457167720e-22 petab = -4.787836794e-28
+ u0 = 1.231769894e-02 lu0 = -3.808197859e-9
+ ua = -2.809317911e-10 lua = -3.619165246e-16
+ ub = 9.337272840e-19 lub = -2.517657501e-25
+ uc = -7.496753916e-11 luc = 1.023045924e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.949154737e+04 lvsat = -1.210264538e-02 wvsat = -4.656612873e-16
+ a0 = 1.349266482e+00 la0 = -2.270095072e-7
+ ags = 1.615750419e-01 lags = 3.344389646e-7
+ a1 = 0.0
+ a2 = 6.001569926e-01 la2 = 3.995391301e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.083405178e-02 lketa = -2.858845418e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.592302506e-01 lpclm = 3.466122321e-7
+ pdiblc1 = 7.407420150e-01 lpdiblc1 = -7.012262346e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.203234000e-01 ldrout = 8.790300377e-7
+ pscbe1 = 7.981743154e+08 lpscbe1 = -1.186332945e+1
+ pscbe2 = 9.526279703e-09 lpscbe2 = -3.492672025e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.883960260e+00 lbeta0 = 1.782957602e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.471808281e-10 lagidl = 7.546826683e-16 pagidl = -1.654361225e-36
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.587827164e-01 lkt1 = -2.026711633e-8
+ kt2 = -5.616202393e-02 lkt2 = 7.597254838e-9
+ at = 9.660944576e+04 lat = -3.482208970e-2
+ ute = 9.121531202e-01 lute = -1.958872090e-06 wute = 1.776356839e-21 pute = 2.664535259e-27
+ ua1 = 6.057818692e-09 lua1 = -6.483453838e-15
+ ub1 = -4.209009179e-18 lub1 = 5.100143366e-24 pub1 = 2.465190329e-44
+ uc1 = -1.262217768e-10 luc1 = 1.929986004e-16 puc1 = 4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.104 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.061395626e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.098818878e-8
+ k1 = 5.226190584e-01 lk1 = -6.426641356e-9
+ k2 = -5.745305410e-03 lk2 = 1.678201184e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.233157705e+00 ldsub = -4.560437967e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.128704363e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.505683220e-9
+ nfactor = {2.446759293e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.834978225e-7
+ eta0 = -1.229902487e-02 leta0 = 2.321282851e-7
+ etab = -1.649900875e+00 letab = 8.234112028e-7
+ u0 = 1.037583596e-02 lu0 = -1.867762149e-9
+ ua = -8.643992354e-11 lua = -5.562654406e-16
+ ub = 1.281983108e-19 lub = 5.531711593e-25
+ uc = -9.823827214e-11 luc = 3.348408823e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.177272666e+04 lvsat = 6.910189940e-2
+ a0 = 1.496294625e+00 la0 = -3.739295848e-7
+ ags = -2.563720021e-01 lags = 7.520788176e-7
+ a1 = 0.0
+ a2 = 1.048426564e+00 la2 = -4.840096337e-8
+ b0 = -8.757847307e-17 lb0 = 8.751410289e-23
+ b1 = -3.641038050e-20 lb1 = 3.638361887e-26
+ keta = 1.074273877e-02 lketa = -2.441977703e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.551875389e+00 lpclm = -7.452298123e-7
+ pdiblc1 = 6.240057999e-02 lpdiblc1 = -2.338338057e-8
+ pdiblc2 = 7.601803479e-04 lpdiblc2 = -3.299376654e-10
+ pdiblcb = -1.455489873e-02 lpdiblcb = -1.043742412e-8
+ drout = 1.037783741e+00 ldrout = -3.775597026e-8
+ pscbe1 = 8.238558016e+08 lpscbe1 = -3.752593977e+1
+ pscbe2 = 3.695351837e-09 lpscbe2 = 5.477374932e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.610435717e+00 lbeta0 = 1.057016105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.015367036e-09 lagidl = -5.069372234e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.243417019e-01 lkt1 = -5.468281666e-8
+ kt2 = -6.234897865e-02 lkt2 = 1.377966215e-8
+ at = 8.491634698e+04 lat = -2.313758535e-2
+ ute = -1.893419934e+00 lute = 8.446388674e-7
+ ua1 = -3.353153283e-09 lua1 = 2.920601073e-15 pua1 = 3.308722450e-36
+ ub1 = 4.101751512e-18 lub1 = -3.204508915e-24
+ uc1 = 3.188735465e-10 luc1 = -2.517695777e-16 wuc1 = 8.271806126e-31 puc1 = 8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.105 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.003044247e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.144612533e-9
+ k1 = 4.418300685e-01 lk1 = 3.390847368e-8
+ k2 = 1.155743619e-02 lk2 = -6.960452102e-09 pk2 = -6.938893904e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.437694134e-01 ldsub = 2.314077213e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.743790865e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.671170052e-8
+ nfactor = {1.493771142e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.922958066e-7
+ eta0 = 4.153918492e-01 leta0 = 1.859720084e-8
+ etab = -1.234637215e-03 letab = 2.898534902e-10
+ u0 = 6.420346145e-03 lu0 = 1.070754753e-10
+ ua = -1.097309096e-09 lua = -5.157384327e-17
+ ub = 8.845879618e-19 lub = 1.755322802e-25
+ uc = -6.126448109e-11 luc = 1.502436844e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.347319152e+05 lvsat = -9.035390602e-3
+ a0 = 8.788192068e-01 la0 = -6.564572002e-08 wa0 = 7.105427358e-21
+ ags = 9.950076829e-01 lags = 1.273087392e-7
+ a1 = 0.0
+ a2 = 1.106485264e+00 la2 = -7.738764019e-8
+ b0 = 1.751569461e-16 lb0 = -4.366049618e-23
+ b1 = 7.282076101e-20 lb1 = -1.815166699e-26
+ keta = -4.464049317e-02 lketa = 3.231132265e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.170588133e-01 lpclm = 2.877166222e-07 wpclm = -1.776356839e-21 ppclm = -6.661338148e-28
+ pdiblc1 = -3.723560082e-01 lpdiblc1 = 1.936753674e-07 wpdiblc1 = -4.440892099e-22 ppdiblc1 = -5.551115123e-29
+ pdiblc2 = -8.352921763e-03 lpdiblc2 = 4.219915260e-09 wpdiblc2 = -1.214306433e-23 ppdiblc2 = 1.062518129e-29
+ pdiblcb = 2.163563710e-01 lpdiblcb = -1.257233392e-07 wpdiblcb = -8.881784197e-22 ppdiblcb = -3.330669074e-28
+ drout = 1.394365649e+00 ldrout = -2.157848363e-7
+ pscbe1 = 6.975643340e+08 lpscbe1 = 2.552696980e+1
+ pscbe2 = 2.047062388e-08 lpscbe2 = -2.897931263e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.545750116e+00 lbeta0 = 9.078136138e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.114932433e-12 lagidl = 5.566467413e-19
+ bgidl = 7.608364006e+08 lbgidl = 1.194060145e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.448437920e-01 lkt1 = 5.479659363e-9
+ kt2 = -1.673808726e-02 lkt2 = -8.992259540e-9
+ at = 9.344592137e+03 lat = 1.459274684e-2
+ ute = 4.294170626e-01 lute = -3.150723455e-07 pute = 4.440892099e-28
+ ua1 = 4.691787198e-09 lua1 = -1.095956137e-15
+ ub1 = -4.457768141e-18 lub1 = 1.068959664e-24 pub1 = -6.162975822e-45
+ uc1 = -2.726704746e-10 luc1 = 4.356764796e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.106 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.370038979e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.953266022e-8
+ k1 = -7.867298771e-01 lk1 = 3.401454685e-7
+ k2 = 5.163552748e-01 lk2 = -1.327888854e-07 wk2 = 1.332267630e-21 pk2 = 3.330669074e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.000619209e+00 ldsub = -3.031133087e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-4.236570348e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.961801644e-8
+ nfactor = {2.329249601e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.065806301e-7
+ eta0 = 1.182779486e+00 leta0 = -1.726856784e-7
+ etab = 6.983305247e-02 letab = -1.742483418e-08 wetab = 3.122502257e-23 petab = 4.987329993e-30
+ u0 = 1.090619245e-02 lu0 = -1.011089003e-9
+ ua = -7.315707161e-10 lua = -1.427396205e-16
+ ub = 1.816775866e-18 lub = -5.682953778e-26
+ uc = -3.744427283e-12 luc = 6.866322317e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.645397497e+05 lvsat = -1.646544047e-2
+ a0 = -7.106838808e-01 la0 = 3.305617671e-7
+ ags = 2.160686824e+00 lags = -1.632542721e-7
+ a1 = 0.0
+ a2 = 1.182249385e+00 la2 = -9.627298368e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.147850760e-01 lketa = 2.071572171e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.759335117e-01 lpclm = -9.654609648e-9
+ pdiblc1 = 1.011312282e+00 lpdiblc1 = -1.512247090e-7
+ pdiblc2 = 2.065758340e-02 lpdiblc2 = -3.011388309e-9
+ pdiblcb = -5.326526217e-02 lpdiblcb = -5.851610281e-8
+ drout = -6.783330112e-01 ldrout = 3.008663952e-7
+ pscbe1 = 7.999049073e+08 lpscbe1 = 1.704680709e-2
+ pscbe2 = 1.260034585e-08 lpscbe2 = -9.361464102e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.034019748e+01 lbeta0 = -3.565115620e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -5.832314471e-10 lagidl = 1.456579198e-16 wagidl = 1.214921525e-30 pagidl = -3.812785636e-37
+ bgidl = 1.854155600e+09 lbgidl = -1.531201959e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.885198056e-01 lkt1 = -8.559939107e-9
+ kt2 = 5.844844661e-02 lkt2 = -2.773363090e-8
+ at = 1.360818822e+05 lat = -1.699842378e-2
+ ute = -2.843863486e+00 lute = 5.008419304e-7
+ ua1 = -8.536520982e-10 lua1 = 2.863277894e-16 pua1 = -8.271806126e-37
+ ub1 = 6.073535279e-19 lub1 = -1.935978887e-25
+ uc1 = -2.923808962e-10 luc1 = 4.848076619e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.107 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-1.827232769e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.401173440e-07 wvth0 = 6.184766960e-07 pvth0 = -1.213853287e-13
+ k1 = 2.281609485e+00 lk1 = -2.298055923e-07 wk1 = -1.014360024e-06 pk1 = 1.990833701e-13
+ k2 = 1.256901662e+00 lk2 = -2.907248142e-07 wk2 = -1.283256875e-06 pk2 = 2.518584105e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.673345986e-01 ldsub = -5.055444706e-08 wdsub = -2.231485290e-07 pdsub = 4.379624604e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {4.226662076e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.455928640e-07 wvoff = -6.426456296e-07 pvoff = 1.261288445e-13
+ nfactor = {2.394425086e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.989599690e-06 wnfactor = -1.761006278e-05 pnfactor = 3.456238971e-12
+ eta0 = 8.493794629e-01 leta0 = -1.236269948e-07 weta0 = -5.456882494e-07 peta0 = 1.070995043e-13
+ etab = -5.930895019e-01 letab = 1.110312348e-07 wetab = 4.900906812e-07 petab = -9.618764755e-14
+ u0 = 9.439774857e-02 lu0 = -1.749344253e-08 wu0 = -7.721590034e-08 pu0 = 1.515477868e-14
+ ua = 9.637465968e-09 lua = -2.191354842e-15 wua = -9.672617624e-15 pua = 1.898396298e-21
+ ub = -3.355017955e-18 lub = 9.528233363e-25 wub = 4.205753125e-24 pub = -8.254421370e-31
+ uc = 2.575474367e-12 luc = -4.886287819e-19 wuc = -2.156797475e-18 puc = 4.233038565e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.541369842e+06 lvsat = 5.130484602e-01 wvsat = 2.264591565e+00 pvsat = -4.444600634e-7
+ a0 = 8.829508915e+00 la0 = -1.510496446e-06 wa0 = -6.667318241e-06 pa0 = 1.308561215e-12
+ ags = 1.249999977e+00 lags = 6.121020135e-15 wags = 6.816088671e-14 pags = -1.337759414e-20
+ a1 = 0.0
+ a2 = -5.130950833e+00 la2 = 1.133657529e-06 wa2 = 5.003954457e-06 pa2 = -9.821011215e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.686950307e-02 lketa = -9.046907693e-09 wketa = -3.993285855e-08 pketa = 7.837422483e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.166966472e-01 lpclm = 1.055950768e-09 wpclm = 4.660894300e-09 ppclm = -9.147704198e-16
+ pdiblc1 = 6.910359467e-01 lpdiblc1 = -1.027065663e-07 wpdiblc1 = -4.533459654e-07 ppdiblc1 = 8.897594590e-14
+ pdiblc2 = 4.055076873e-02 lpdiblc2 = -7.201299321e-09 wpdiblc2 = -3.178648372e-08 ppdiblc2 = 6.238574228e-15
+ pdiblcb = -1.890403849e+00 lpdiblcb = 2.965007219e-07 wpdiblcb = 1.308751058e-06 ppdiblcb = -2.568620264e-13
+ drout = 1.000002350e+00 ldrout = -4.306521504e-13 wdrout = -1.152224826e-12 pdrout = 2.261414096e-19
+ pscbe1 = 8.000000125e+08 lpscbe1 = -2.447006226e-06 wpscbe1 = -1.052743530e-05 ppscbe1 = 2.066169739e-12
+ pscbe2 = -2.698060633e-08 lpscbe2 = 6.743432838e-15 wpscbe2 = 2.976545202e-14 ppscbe2 = -5.841916441e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.272015552e+01 lbeta0 = -8.574226144e-07 wbeta0 = -3.784657842e-06 pbeta0 = 7.427958714e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 5.662539482e-08 lagidl = -1.106858013e-14 wagidl = -4.885661624e-14 pagidl = 9.588843786e-21
+ bgidl = 1.000000294e+09 lbgidl = -4.915885162e-05 wbgidl = -7.498443604e-06 pbgidl = 1.471687317e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 5.380173401e-01 lkt1 = -2.108450054e-07 wkt1 = -9.306680303e-07 pkt1 = 1.826575610e-13
+ kt2 = -9.625899335e-02 lkt2 = -1.839462804e-15 wkt2 = -2.120583531e-14 pkt2 = 4.161963219e-21
+ at = 7.216409615e+05 lat = -1.335351655e-01 wat = -5.894230514e-01 pat = 1.156831152e-7
+ ute = -1.661431450e+00 lute = 3.162675854e-07 wute = 1.396002169e-06 pute = -2.739863657e-13
+ ua1 = 7.435796699e-10 lua1 = 3.992814052e-23 wua1 = -4.319688036e-22 pua1 = 8.478034825e-29
+ ub1 = -4.726028342e-19 lub1 = 5.349365731e-31 wub1 = 1.839635587e-30 pub1 = -3.610560804e-37
+ uc1 = -2.193903888e-11 luc1 = 7.270256460e-24 wuc1 = 2.325127940e-23 puc1 = -4.563412337e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.108 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.109 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.124648838e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.706194604e-7
+ k1 = 4.210818616e-01 lk1 = 2.114671972e-7
+ k2 = 2.113420949e-02 lk2 = 8.596014224e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = -6.776263578e-27 pcit = 3.794707604e-31
+ voff = {-2.804004741e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.598181832e-7
+ nfactor = {1.983803335e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.424216791e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.153077275e-02 lu0 = -2.044270362e-8
+ ua = -9.098047201e-10 lua = 1.854443048e-15
+ ub = 1.491779338e-18 lub = -5.043522411e-24
+ uc = -1.282516351e-10 luc = 4.517563002e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.672490943e+04 lvsat = 1.068582539e+0
+ a0 = 1.566615238e+00 la0 = -2.052229338e-6
+ ags = 6.394720045e-02 lags = 9.868197240e-7
+ a1 = 0.0
+ a2 = 1.083322921e+00 la2 = -2.266375124e-6
+ b0 = -2.161420565e-07 lb0 = 1.728977587e-12
+ b1 = 9.955134135e-10 lb1 = -7.963375606e-15
+ keta = 4.018068624e-02 lketa = -3.363761825e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.896493835e-02 lpclm = 1.679237053e-06 wpclm = -1.110223025e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.915673984e-03 lpdiblc2 = -1.276983438e-8
+ pdiblcb = -2.715826998e-01 lpdiblcb = 9.316197581e-07 wpdiblcb = -1.776356839e-21
+ drout = 0.56
+ pscbe1 = 8.000324970e+08 lpscbe1 = -6.499163959e-1
+ pscbe2 = 1.315044923e-08 lpscbe2 = -6.179421357e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.666054167e-11 lalpha0 = 1.333161838e-15
+ alpha1 = -6.666054167e-11 lalpha1 = 1.333161838e-15
+ beta0 = 4.581282086e+01 lbeta0 = -3.162447948e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.870274718e-09 lagidl = -1.939963340e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.235849912e-01 legidl = 1.047131499e-5
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365691544e-01 lkt1 = -3.361567574e-08 wkt1 = 3.552713679e-21
+ kt2 = -6.267063968e-02 lkt2 = 8.248976200e-08 wkt2 = 4.440892099e-22
+ at = 1.183123185e+05 lat = -9.464115887e-1
+ ute = -5.012560544e-02 lute = -6.570637432e-7
+ ua1 = 2.268500750e-09 lua1 = -3.565883958e-15
+ ub1 = -1.570875991e-18 lub1 = 6.839268476e-24
+ uc1 = -4.380619758e-11 luc1 = 2.803336491e-16 wuc1 = 2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.110 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.069866256e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.239906809e-8
+ k1 = 4.556237202e-01 lk1 = -6.484228401e-8
+ k2 = 2.007683582e-02 lk2 = 1.705422642e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.164179846e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.199470589e-8
+ nfactor = {2.378038919e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.167837078e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.443397737e-03 lu0 = 4.254027232e-9
+ ua = -7.572954228e-10 lua = 6.344807637e-16
+ ub = 8.922232633e-19 lub = -2.475144842e-25
+ uc = -7.084368051e-11 luc = -7.465141979e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.671623623e+05 lvsat = -8.547403617e-1
+ a0 = 1.370094967e+00 la0 = -4.802116133e-7
+ ags = 1.321801322e-01 lags = 4.410064215e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.426888399e-04 lketa = -8.219334060e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.401119263e-01 lpclm = -7.931506930e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.387319811e-03 lpdiblc2 = 1.365168829e-08 wpdiblc2 = 3.469446952e-24 ppdiblc2 = -1.387778781e-29
+ pdiblcb = -2.488330300e-01 lpdiblcb = 7.496391204e-07 wpdiblcb = -1.776356839e-21
+ drout = 0.56
+ pscbe1 = 1.224636900e+09 lpscbe1 = -3.397173053e+3
+ pscbe2 = -1.698011262e-08 lpscbe2 = 1.792281353e-13 ppscbe2 = 2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.446751046e+00 lbeta0 = 2.265262463e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.904539975e-10 lagidl = -1.962669803e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.670754974e+00 legidl = -6.281865390e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.063193317e-01 lkt1 = -2.755920237e-7
+ kt2 = -4.841666844e-02 lkt2 = -3.153153126e-8
+ at = -9.065933829e+04 lat = 7.252080717e-1
+ ute = -1.645263111e-01 lute = 2.580578176e-7
+ ua1 = 5.778773827e-10 lua1 = 9.957860376e-15
+ ub1 = 8.146409535e-19 lub1 = -1.224311373e-23 pub1 = 4.930380658e-44
+ uc1 = -1.163111597e-11 luc1 = 2.295664482e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.111 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063199473e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.736836213e-9
+ k1 = 4.427665361e-01 lk1 = -1.342299740e-8
+ k2 = 2.238297990e-02 lk2 = 7.831345119e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.585912374e-01 ldsub = -1.194145485e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.482687602e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.538498620e-8
+ nfactor = {9.059919706e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.719268760e-6
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394757071e-01 letab = 2.778517638e-7
+ u0 = 8.601632882e-03 lu0 = 3.621202956e-9
+ ua = -7.352853466e-10 lua = 5.464566366e-16
+ ub = 8.528601283e-19 lub = -9.009087610e-26
+ uc = -7.556913799e-11 luc = 1.143321474e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.264314745e+00 la0 = -5.716847236e-8
+ ags = 1.560797535e-01 lags = 3.454255025e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.464757958e-03 lketa = -3.744375028e-08 pketa = 5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.488073345e-01 lpclm = 2.361946495e-06 wpclm = 1.776356839e-21 ppclm = -4.440892099e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.621872386e-03 lpdiblc2 = -6.381398745e-9
+ pdiblcb = -9.776424111e-02 lpdiblcb = 1.454750005e-7
+ drout = 0.56
+ pscbe1 = -4.171210305e+07 lpscbe1 = 1.667292191e+3
+ pscbe2 = 4.631193739e-08 lpscbe2 = -7.389354511e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.144527102e+01 lbeta0 = -9.335576356e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.690680066e-10 lagidl = -2.774355581e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815376811e-01 lkt1 = 2.522608815e-8
+ kt2 = -6.023855242e-02 lkt2 = 1.574731557e-8
+ at = 1.021557796e+05 lat = -4.591068088e-2
+ ute = -1.323451088e-01 lute = 1.293566616e-7
+ ua1 = 3.320607059e-09 lua1 = -1.011042424e-15
+ ub1 = -2.835183653e-18 lub1 = 2.353502076e-24
+ uc1 = 1.789645493e-11 luc1 = -9.513193603e-17 wuc1 = 5.169878828e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.112 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.080253346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.983204748e-8
+ k1 = 3.559763493e-01 lk1 = 1.600935854e-7
+ k2 = 5.664373486e-02 lk2 = -6.066498314e-08 wk2 = -2.220446049e-22 pk2 = 2.220446049e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.538016126e-01 ldsub = 1.029822606e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.107617634e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.985602103e-10
+ nfactor = {2.269123695e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.992787282e-9
+ eta0 = -2.188386675e-01 leta0 = 4.385161211e-07 weta0 = 3.608224830e-22 peta0 = 4.163336342e-29
+ etab = 8.242798594e-01 letab = -1.648951009e-06 wetab = -1.679212325e-21 petab = -9.228728892e-28
+ u0 = 1.231769894e-02 lu0 = -3.808197859e-9
+ ua = -2.809317911e-10 lua = -3.619165246e-16
+ ub = 9.337272840e-19 lub = -2.517657501e-25
+ uc = -7.496753916e-11 luc = 1.023045924e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.949154737e+04 lvsat = -1.210264538e-02 wvsat = -4.656612873e-16
+ a0 = 1.349266482e+00 la0 = -2.270095072e-7
+ ags = 1.615750419e-01 lags = 3.344389646e-7
+ a1 = 0.0
+ a2 = 6.001569926e-01 la2 = 3.995391301e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.083405178e-02 lketa = -2.858845418e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.592302506e-01 lpclm = 3.466122321e-7
+ pdiblc1 = 7.407420150e-01 lpdiblc1 = -7.012262346e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.203234000e-01 ldrout = 8.790300377e-7
+ pscbe1 = 7.981743154e+08 lpscbe1 = -1.186332945e+1
+ pscbe2 = 9.526279703e-09 lpscbe2 = -3.492672025e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.883960260e+00 lbeta0 = 1.782957602e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.471808281e-10 lagidl = 7.546826683e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.587827164e-01 lkt1 = -2.026711633e-8
+ kt2 = -5.616202393e-02 lkt2 = 7.597254838e-9
+ at = 9.660944576e+04 lat = -3.482208970e-2
+ ute = 9.121531202e-01 lute = -1.958872090e-06 pute = -2.664535259e-27
+ ua1 = 6.057818692e-09 lua1 = -6.483453838e-15
+ ub1 = -4.209009179e-18 lub1 = 5.100143366e-24 wub1 = 2.465190329e-38
+ uc1 = -1.262217768e-10 luc1 = 1.929986004e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.113 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.061395626e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.098818878e-8
+ k1 = 5.226190584e-01 lk1 = -6.426641356e-9
+ k2 = -5.745305410e-03 lk2 = 1.678201184e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.233157705e+00 ldsub = -4.560437967e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.128704363e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.505683220e-9
+ nfactor = {2.446759293e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.834978225e-7
+ eta0 = -1.229902487e-02 leta0 = 2.321282851e-7
+ etab = -1.649900875e+00 letab = 8.234112028e-7
+ u0 = 1.037583596e-02 lu0 = -1.867762149e-9
+ ua = -8.643992354e-11 lua = -5.562654406e-16
+ ub = 1.281983108e-19 lub = 5.531711593e-25
+ uc = -9.823827214e-11 luc = 3.348408823e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.177272666e+04 lvsat = 6.910189940e-02 pvsat = 2.328306437e-22
+ a0 = 1.496294625e+00 la0 = -3.739295848e-7
+ ags = -2.563720021e-01 lags = 7.520788176e-7
+ a1 = 0.0
+ a2 = 1.048426564e+00 la2 = -4.840096337e-8
+ b0 = -8.757847307e-17 lb0 = 8.751410289e-23
+ b1 = -3.641038050e-20 lb1 = 3.638361887e-26
+ keta = 1.074273877e-02 lketa = -2.441977703e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.551875389e+00 lpclm = -7.452298123e-7
+ pdiblc1 = 6.240057999e-02 lpdiblc1 = -2.338338057e-8
+ pdiblc2 = 7.601803479e-04 lpdiblc2 = -3.299376654e-10
+ pdiblcb = -1.455489873e-02 lpdiblcb = -1.043742412e-8
+ drout = 1.037783741e+00 ldrout = -3.775597026e-8
+ pscbe1 = 8.238558016e+08 lpscbe1 = -3.752593977e+1
+ pscbe2 = 3.695351837e-09 lpscbe2 = 5.477374932e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.610435717e+00 lbeta0 = 1.057016105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.015367036e-09 lagidl = -5.069372234e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.243417019e-01 lkt1 = -5.468281666e-8
+ kt2 = -6.234897865e-02 lkt2 = 1.377966215e-8
+ at = 8.491634698e+04 lat = -2.313758535e-2
+ ute = -1.893419934e+00 lute = 8.446388674e-7
+ ua1 = -3.353153283e-09 lua1 = 2.920601073e-15 pua1 = 3.308722450e-36
+ ub1 = 4.101751512e-18 lub1 = -3.204508915e-24
+ uc1 = 3.188735465e-10 luc1 = -2.517695777e-16 puc1 = 8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.114 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.003044247e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.144612533e-9
+ k1 = 4.418300685e-01 lk1 = 3.390847368e-8
+ k2 = 1.155743619e-02 lk2 = -6.960452102e-09 pk2 = 2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.437694134e-01 ldsub = 2.314077213e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.743790865e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.671170052e-8
+ nfactor = {1.493771142e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.922958066e-7
+ eta0 = 4.153918492e-01 leta0 = 1.859720084e-8
+ etab = -1.234637215e-03 letab = 2.898534902e-10
+ u0 = 6.420346145e-03 lu0 = 1.070754753e-10
+ ua = -1.097309096e-09 lua = -5.157384327e-17
+ ub = 8.845879618e-19 lub = 1.755322802e-25
+ uc = -6.126448109e-11 luc = 1.502436844e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.347319152e+05 lvsat = -9.035390602e-3
+ a0 = 8.788192068e-01 la0 = -6.564572002e-8
+ ags = 9.950076829e-01 lags = 1.273087392e-7
+ a1 = 0.0
+ a2 = 1.106485264e+00 la2 = -7.738764019e-8
+ b0 = 1.751569461e-16 lb0 = -4.366049618e-23
+ b1 = 7.282076101e-20 lb1 = -1.815166699e-26
+ keta = -4.464049317e-02 lketa = 3.231132265e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.170588133e-01 lpclm = 2.877166222e-07 wpclm = 1.776356839e-21 ppclm = -8.881784197e-28
+ pdiblc1 = -3.723560082e-01 lpdiblc1 = 1.936753674e-07 wpdiblc1 = 2.220446049e-22 ppdiblc1 = 2.220446049e-28
+ pdiblc2 = -8.352921763e-03 lpdiblc2 = 4.219915260e-09 wpdiblc2 = -6.071532166e-24 ppdiblc2 = 5.421010862e-30
+ pdiblcb = 2.163563710e-01 lpdiblcb = -1.257233392e-07 ppdiblcb = -4.440892099e-28
+ drout = 1.394365649e+00 ldrout = -2.157848363e-7
+ pscbe1 = 6.975643340e+08 lpscbe1 = 2.552696980e+1
+ pscbe2 = 2.047062388e-08 lpscbe2 = -2.897931263e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.545750116e+00 lbeta0 = 9.078136138e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.114932433e-12 lagidl = 5.566467413e-19
+ bgidl = 7.608364006e+08 lbgidl = 1.194060145e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.448437920e-01 lkt1 = 5.479659363e-9
+ kt2 = -1.673808726e-02 lkt2 = -8.992259540e-9
+ at = 9.344592137e+03 lat = 1.459274684e-2
+ ute = 4.294170626e-01 lute = -3.150723455e-07 pute = 4.440892099e-28
+ ua1 = 4.691787198e-09 lua1 = -1.095956137e-15
+ ub1 = -4.457768141e-18 lub1 = 1.068959664e-24
+ uc1 = -2.726704746e-10 luc1 = 4.356764796e-17 wuc1 = 1.654361225e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.115 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {1.251447606e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.701105243e-07 wvth0 = -1.809250599e-06 pvth0 = 4.509828506e-13
+ k1 = -1.114561074e+00 lk1 = 4.218623118e-07 wk1 = 2.840040997e-07 pk1 = -7.079228191e-14
+ k2 = -9.317975967e-01 lk2 = 2.281849402e-07 wk2 = 1.254552210e-06 pk2 = -3.127159567e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.044442743e+00 ldsub = -5.633019819e-07 wdsub = -9.042768531e-07 pdsub = 2.254045698e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-4.514098852e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.234238151e-08 wvoff = 3.543598831e-07 pvoff = -8.832951627e-14
+ nfactor = {-2.480166249e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.282859310e-06 wnfactor = 2.350383472e-06 pnfactor = -5.858683361e-13
+ eta0 = 3.490815564e+00 leta0 = -7.479982914e-07 weta0 = -1.999479351e-06 peta0 = 4.984002204e-13
+ etab = 2.926356743e-01 letab = -7.296172971e-08 wetab = -1.930165849e-07 petab = 4.811227904e-14
+ u0 = -1.891672623e-02 lu0 = 6.422720822e-09 wu0 = 2.583595233e-08 pu0 = -6.439998657e-15
+ ua = -7.260372955e-09 lua = 1.484662270e-15 wua = 5.655979725e-15 pua = -1.409837786e-21
+ ub = 7.146304487e-18 lub = -1.385294490e-24 wub = -4.617034599e-24 pub = 1.150865129e-30
+ uc = -1.164889050e-10 luc = 2.878988446e-17 wuc = 9.767189395e-17 puc = -2.434618465e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.204121918e+05 lvsat = -1.051719848e-01 wvsat = -3.082965671e-01 pvsat = 7.684754379e-8
+ a0 = -2.896295838e+00 la0 = 8.753583316e-07 wa0 = 1.893421866e-06 pa0 = -4.719638013e-13
+ ags = 2.160686853e+00 lags = -1.632542791e-07 wags = -2.456459924e-14 pags = 6.123094920e-21
+ a1 = 0.0
+ a2 = 2.051783901e+00 la2 = -3.130175048e-07 wa2 = -7.532881856e-07 pa2 = 1.877683796e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.285162498e-01 lketa = 4.906492273e-08 wketa = 9.852668060e-08 pketa = -2.455925304e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.649693630e-01 lpclm = -6.921631119e-09 wpclm = 9.498373599e-09 ppclm = -2.367612095e-15
+ pdiblc1 = 2.585423770e+00 lpdiblc1 = -5.435956090e-07 wpdiblc1 = -1.363671671e-06 ppdiblc1 = 3.399156191e-13
+ pdiblc2 = -1.372744820e-03 lpdiblc2 = 2.480001454e-09 wpdiblc2 = 1.908513770e-08 ppdiblc2 = -4.757256849e-15
+ pdiblcb = -6.433784370e+00 lpdiblcb = 1.531923993e-06 wpdiblcb = 5.527520270e-06 ppdiblcb = -1.377817340e-12
+ drout = -6.783342909e-01 ldrout = 3.008667142e-07 wdrout = 1.108640078e-12 pdrout = -2.763451690e-19
+ pscbe1 = 7.999049111e+08 lpscbe1 = 1.704585167e-02 wpscbe1 = -3.320541382e-06 ppscbe1 = 8.276977539e-13
+ pscbe2 = -6.083460749e-09 lpscbe2 = 3.721072641e-15 wpscbe2 = 1.618600586e-14 ppscbe2 = -4.034604751e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.036110947e+01 lbeta0 = -3.617241888e-07 wbeta0 = -1.811630667e-08 pbeta0 = 4.515761183e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.532708909e-08 lagidl = 6.313435594e-15 wagidl = 2.143590080e-14 pagidl = -5.343219813e-21
+ bgidl = 1.854155615e+09 lbgidl = -1.531201994e+02 wbgidl = -1.232455444e-05 pbgidl = 3.072078705e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.186979074e-01 lkt1 = 9.866840543e-08 wkt1 = 3.726684517e-07 pkt1 = -9.289320161e-14
+ kt2 = 4.405273520e-01 lkt2 = -1.229725292e-07 wkt2 = -3.309995407e-07 pkt2 = 8.250660050e-14
+ at = -5.699521945e+04 lat = 3.112893997e-02 wat = 1.672650101e-01 pat = -4.169331274e-8
+ ute = -6.484173388e+00 lute = 1.408243778e-06 wute = 3.153644153e-06 pute = -7.860931097e-13
+ ua1 = -4.160807027e-09 lua1 = 1.110685763e-15 wua1 = 2.865028001e-15 pua1 = -7.141512047e-22
+ ub1 = 3.621521657e-18 lub1 = -9.449245073e-25 wub1 = -2.611210020e-24 pub1 = 6.508832657e-31
+ uc1 = -3.542388178e-10 luc1 = 6.389978101e-17 wuc1 = 5.358825975e-17 puc1 = -1.335767757e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.116 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-5.146198521e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.314589576e-07 wvth0 = 3.493736555e-06 pvth0 = -5.470404647e-13
+ k1 = 1.238729295e+00 lk1 = -3.133406210e-13 wk1 = -1.109004007e-07 pk1 = 2.992794492e-19
+ k2 = 1.864770599e+00 lk2 = -2.990443570e-07 wk2 = -1.809861030e-06 pk2 = 2.590657303e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -9.785075347e-02 ldsub = 1.381405950e-12 wdsub = 3.531095238e-07 pdsub = -8.748370881e-19
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.594266927e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.590003684e-14 wvoff = -1.383715650e-07 pvoff = -1.447315334e-20
+ nfactor = {4.676024599e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.209075454e-12 wnfactor = -9.177671528e-07 pnfactor = -3.628686926e-18
+ eta0 = -6.817674743e-01 leta0 = -2.113539139e-13 weta0 = 7.807627161e-07 peta0 = 1.382324175e-19
+ etab = -1.143701283e-01 letab = 1.811845247e-13 wetab = 7.537034328e-08 petab = -1.134735428e-19
+ u0 = -1.317756369e-02 lu0 = 5.905401450e-09 wu0 = 1.597788358e-08 pu0 = -5.115920646e-15
+ ua = 1.021738640e-09 lua = -3.335463627e-20 wua = -2.208709651e-15 pua = 2.819723014e-26
+ ub = -5.813339295e-19 lub = 6.692371254e-31 wub = 1.802877370e-24 pub = -4.266986107e-37
+ uc = 4.411068443e-11 luc = -1.020136723e-24 wuc = -3.813924838e-17 puc = -2.370290690e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.122374658e+05 lvsat = -1.135412075e-01 wvsat = -3.807850891e-01 pvsat = 9.836208476e-8
+ a0 = 1.986741243e+00 la0 = 7.547192808e-13 wa0 = -7.393464937e-07 pa0 = -6.365323699e-19
+ ags = 1.249999986e+00 lags = 2.225164053e-15 wags = 6.055660151e-14 pags = -1.000255878e-20
+ a1 = 0.0
+ a2 = 3.056678521e-01 la2 = -1.244513470e-14 wa2 = 2.941464508e-07 pa2 = 1.039600406e-20
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.518476887e-02 lketa = -9.894333676e-14 wketa = -3.847335310e-08 pketa = 6.350102641e-20
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.263578362e-01 lpclm = 7.031776406e-14 wpclm = -3.708709670e-09 ppclm = -4.851528956e-20
+ pdiblc1 = -4.469354772e-01 lpdiblc1 = 2.972046333e-13 wpdiblc1 = 5.324923348e-07 ppdiblc1 = -2.424055117e-19
+ pdiblc2 = 1.246149974e-02 lpdiblc2 = 6.133613645e-15 wpdiblc2 = -7.452412935e-09 ppdiblc2 = -3.102969909e-21
+ pdiblcb = 2.111796305e+00 lpdiblcb = 5.176975861e-13 wpdiblcb = -2.158402962e-06 ppdiblcb = -3.415426342e-19
+ drout = 1.000004188e+00 ldrout = -6.933270242e-13 wdrout = -2.744574942e-12 pdrout = 4.536998048e-19
+ pscbe1 = 7.999999861e+08 lpscbe1 = 2.439033508e-06 wpscbe1 = 1.233615112e-05 ppscbe1 = -2.166675568e-12
+ pscbe2 = 1.467392486e-08 lpscbe2 = -9.850363196e-23 wpscbe2 = -6.320368201e-15 ppscbe2 = 4.327755496e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.343284779e+00 lbeta0 = 1.264576326e-12 wbeta0 = 7.077805691e-09 pbeta0 = -7.240887498e-19
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 9.891362726e-09 lagidl = -1.860982455e-22 wagidl = -8.370363432e-15 pagidl = 1.584177415e-28
+ bgidl = 1.000000314e+09 lbgidl = -5.408121490e-05 wbgidl = -2.441311646e-05 pbgidl = 5.735961914e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.682918657e-01 lkt1 = -1.462992962e-13 wkt1 = -1.455214897e-07 pkt1 = 1.294359464e-19
+ kt2 = -2.454538498e-01 lkt2 = -1.194574653e-13 wkt2 = 1.292492733e-07 pkt2 = 1.060558503e-19
+ at = 1.166522731e+05 lat = 2.433537319e-08 wat = -6.531409069e-02 pat = -2.215757710e-14
+ ute = 1.371480169e+00 lute = 4.744966153e-14 wute = -1.231445561e-06 pute = -2.323446102e-21
+ ua1 = 2.034962688e-09 lua1 = 1.209538141e-21 wua1 = -1.118741037e-15 pua1 = -9.284668272e-28
+ ub1 = -1.649583075e-18 lub1 = 9.025072579e-32 wub1 = 1.019633946e-24 pub1 = 2.418060820e-38
+ uc1 = 2.215392550e-12 luc1 = 1.861136381e-23 wuc1 = -2.092525055e-17 puc1 = -1.438834994e-29
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.117 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.118 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.124648838e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.706194604e-7
+ k1 = 4.210818616e-01 lk1 = 2.114671972e-7
+ k2 = 2.113420949e-02 lk2 = 8.596014224e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = 3.388131789e-27 pcit = -1.084202172e-31
+ voff = {-2.804004741e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.598181832e-7
+ nfactor = {1.983803335e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.424216791e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.153077275e-02 lu0 = -2.044270362e-08 wu0 = -5.551115123e-23
+ ua = -9.098047201e-10 lua = 1.854443048e-15
+ ub = 1.491779338e-18 lub = -5.043522411e-24
+ uc = -1.282516351e-10 luc = 4.517563002e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.672490943e+04 lvsat = 1.068582539e+0
+ a0 = 1.566615238e+00 la0 = -2.052229338e-6
+ ags = 6.394720045e-02 lags = 9.868197240e-7
+ a1 = 0.0
+ a2 = 1.083322921e+00 la2 = -2.266375124e-6
+ b0 = -2.161420565e-07 lb0 = 1.728977587e-12
+ b1 = 9.955134135e-10 lb1 = -7.963375606e-15
+ keta = 4.018068624e-02 lketa = -3.363761825e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.896493835e-02 lpclm = 1.679237053e-06 wpclm = -1.110223025e-22 ppclm = 1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.915673984e-03 lpdiblc2 = -1.276983438e-8
+ pdiblcb = -2.715826998e-01 lpdiblcb = 9.316197581e-7
+ drout = 0.56
+ pscbe1 = 8.000324970e+08 lpscbe1 = -6.499163959e-1
+ pscbe2 = 1.315044923e-08 lpscbe2 = -6.179421357e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.666054167e-11 lalpha0 = 1.333161838e-15
+ alpha1 = -6.666054167e-11 lalpha1 = 1.333161838e-15
+ beta0 = 4.581282086e+01 lbeta0 = -3.162447948e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.870274718e-09 lagidl = -1.939963340e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.235849912e-01 legidl = 1.047131499e-05 wegidl = 8.881784197e-22 pegidl = -3.552713679e-27
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365691544e-01 lkt1 = -3.361567574e-8
+ kt2 = -6.267063968e-02 lkt2 = 8.248976200e-8
+ at = 1.183123185e+05 lat = -9.464115887e-1
+ ute = -5.012560544e-02 lute = -6.570637432e-7
+ ua1 = 2.268500750e-09 lua1 = -3.565883958e-15
+ ub1 = -1.570875991e-18 lub1 = 6.839268476e-24
+ uc1 = -4.380619758e-11 luc1 = 2.803336491e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.119 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.069866256e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.239906809e-8
+ k1 = 4.556237202e-01 lk1 = -6.484228401e-8
+ k2 = 2.007683582e-02 lk2 = 1.705422642e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.164179846e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.199470589e-8
+ nfactor = {2.378038919e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.167837078e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.443397737e-03 lu0 = 4.254027232e-9
+ ua = -7.572954228e-10 lua = 6.344807637e-16
+ ub = 8.922232633e-19 lub = -2.475144842e-25
+ uc = -7.084368051e-11 luc = -7.465141979e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.671623623e+05 lvsat = -8.547403617e-1
+ a0 = 1.370094967e+00 la0 = -4.802116133e-7
+ ags = 1.321801322e-01 lags = 4.410064215e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.426888399e-04 lketa = -8.219334060e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.401119263e-01 lpclm = -7.931506930e-07 wpclm = -8.881784197e-22
+ pdiblc1 = 0.39
+ pdiblc2 = -1.387319811e-03 lpdiblc2 = 1.365168829e-08 wpdiblc2 = 1.734723476e-24 ppdiblc2 = 2.775557562e-29
+ pdiblcb = -2.488330300e-01 lpdiblcb = 7.496391204e-7
+ drout = 0.56
+ pscbe1 = 1.224636900e+09 lpscbe1 = -3.397173053e+3
+ pscbe2 = -1.698011262e-08 lpscbe2 = 1.792281353e-13 ppscbe2 = -4.235164736e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.446751046e+00 lbeta0 = 2.265262463e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.904539975e-10 lagidl = -1.962669803e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.670754974e+00 legidl = -6.281865390e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.063193317e-01 lkt1 = -2.755920237e-7
+ kt2 = -4.841666844e-02 lkt2 = -3.153153126e-8
+ at = -9.065933828e+04 lat = 7.252080717e-1
+ ute = -1.645263111e-01 lute = 2.580578176e-7
+ ua1 = 5.778773827e-10 lua1 = 9.957860376e-15
+ ub1 = 8.146409535e-19 lub1 = -1.224311373e-23 pub1 = 2.465190329e-44
+ uc1 = -1.163111597e-11 luc1 = 2.295664482e-17 wuc1 = -5.169878828e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.120 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063199473e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.736836213e-9
+ k1 = 4.427665361e-01 lk1 = -1.342299740e-8
+ k2 = 2.238297990e-02 lk2 = 7.831345119e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.585912374e-01 ldsub = -1.194145485e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.482687602e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.538498620e-8
+ nfactor = {9.059919706e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.719268760e-6
+ eta0 = 1.594707837e-01 leta0 = -3.178247240e-7
+ etab = -1.394757071e-01 letab = 2.778517638e-7
+ u0 = 8.601632881e-03 lu0 = 3.621202956e-9
+ ua = -7.352853466e-10 lua = 5.464566366e-16 wua = -3.308722450e-30
+ ub = 8.528601283e-19 lub = -9.009087610e-26
+ uc = -7.556913799e-11 luc = 1.143321474e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.264314745e+00 la0 = -5.716847236e-8
+ ags = 1.560797535e-01 lags = 3.454255025e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.464757958e-03 lketa = -3.744375028e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.488073345e-01 lpclm = 2.361946495e-06 wpclm = 4.440892099e-22 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 3.621872386e-03 lpdiblc2 = -6.381398745e-9
+ pdiblcb = -9.776424111e-02 lpdiblcb = 1.454750005e-7
+ drout = 0.56
+ pscbe1 = -4.171210305e+07 lpscbe1 = 1.667292191e+3
+ pscbe2 = 4.631193739e-08 lpscbe2 = -7.389354511e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.144527102e+01 lbeta0 = -9.335576356e-06 wbeta0 = 5.684341886e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.690680066e-10 lagidl = -2.774355581e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815376811e-01 lkt1 = 2.522608815e-8
+ kt2 = -6.023855242e-02 lkt2 = 1.574731557e-8
+ at = 1.021557796e+05 lat = -4.591068088e-02 wat = -4.656612873e-16
+ ute = -1.323451088e-01 lute = 1.293566616e-7
+ ua1 = 3.320607059e-09 lua1 = -1.011042424e-15
+ ub1 = -2.835183653e-18 lub1 = 2.353502076e-24
+ uc1 = 1.789645493e-11 luc1 = -9.513193603e-17 puc1 = 1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.121 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.080253346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.983204748e-8
+ k1 = 3.559763493e-01 lk1 = 1.600935854e-7
+ k2 = 5.664373486e-02 lk2 = -6.066498314e-08 pk2 = -2.220446049e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.538016126e-01 ldsub = 1.029822606e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.107617634e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.985602103e-10
+ nfactor = {2.269123695e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.992787282e-9
+ eta0 = -2.188386675e-01 leta0 = 4.385161211e-07 weta0 = 3.295974604e-22 peta0 = -7.285838599e-29
+ etab = 8.242798594e-01 letab = -1.648951009e-06 wetab = 1.477984402e-21 petab = -3.268219029e-27
+ u0 = 1.231769894e-02 lu0 = -3.808197859e-9
+ ua = -2.809317911e-10 lua = -3.619165246e-16
+ ub = 9.337272840e-19 lub = -2.517657501e-25
+ uc = -7.496753916e-11 luc = 1.023045924e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.949154737e+04 lvsat = -1.210264538e-2
+ a0 = 1.349266482e+00 la0 = -2.270095072e-7
+ ags = 1.615750419e-01 lags = 3.344389646e-7
+ a1 = 0.0
+ a2 = 6.001569926e-01 la2 = 3.995391301e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.083405178e-02 lketa = -2.858845418e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.592302506e-01 lpclm = 3.466122321e-7
+ pdiblc1 = 7.407420150e-01 lpdiblc1 = -7.012262346e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.203234000e-01 ldrout = 8.790300377e-7
+ pscbe1 = 7.981743154e+08 lpscbe1 = -1.186332945e+1
+ pscbe2 = 9.526279703e-09 lpscbe2 = -3.492672025e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.883960260e+00 lbeta0 = 1.782957602e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.471808281e-10 lagidl = 7.546826683e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.587827164e-01 lkt1 = -2.026711633e-8
+ kt2 = -5.616202393e-02 lkt2 = 7.597254838e-9
+ at = 9.660944576e+04 lat = -3.482208970e-2
+ ute = 9.121531202e-01 lute = -1.958872090e-06 pute = 1.776356839e-27
+ ua1 = 6.057818692e-09 lua1 = -6.483453838e-15 pua1 = 2.646977960e-35
+ ub1 = -4.209009179e-18 lub1 = 5.100143366e-24
+ uc1 = -1.262217768e-10 luc1 = 1.929986004e-16 wuc1 = 2.067951531e-31 puc1 = 4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.122 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.061395626e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.098818878e-8
+ k1 = 5.226190584e-01 lk1 = -6.426641356e-9
+ k2 = -5.745305410e-03 lk2 = 1.678201184e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.233157705e+00 ldsub = -4.560437967e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.128704363e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.505683220e-9
+ nfactor = {2.446759293e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.834978225e-7
+ eta0 = -1.229902487e-02 leta0 = 2.321282851e-7
+ etab = -1.649900875e+00 letab = 8.234112028e-7
+ u0 = 1.037583596e-02 lu0 = -1.867762149e-9
+ ua = -8.643992354e-11 lua = -5.562654406e-16
+ ub = 1.281983108e-19 lub = 5.531711593e-25
+ uc = -9.823827214e-11 luc = 3.348408823e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.177272666e+04 lvsat = 6.910189940e-2
+ a0 = 1.496294625e+00 la0 = -3.739295848e-7
+ ags = -2.563720021e-01 lags = 7.520788176e-07 pags = 1.776356839e-27
+ a1 = 0.0
+ a2 = 1.048426564e+00 la2 = -4.840096337e-8
+ b0 = -8.757847307e-17 lb0 = 8.751410289e-23
+ b1 = -3.641038050e-20 lb1 = 3.638361887e-26
+ keta = 1.074273877e-02 lketa = -2.441977703e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.551875389e+00 lpclm = -7.452298123e-7
+ pdiblc1 = 6.240057999e-02 lpdiblc1 = -2.338338057e-8
+ pdiblc2 = 7.601803479e-04 lpdiblc2 = -3.299376654e-10
+ pdiblcb = -1.455489873e-02 lpdiblcb = -1.043742412e-8
+ drout = 1.037783741e+00 ldrout = -3.775597026e-8
+ pscbe1 = 8.238558016e+08 lpscbe1 = -3.752593977e+1
+ pscbe2 = 3.695351837e-09 lpscbe2 = 5.477374932e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.610435717e+00 lbeta0 = 1.057016105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.015367036e-09 lagidl = -5.069372234e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.243417019e-01 lkt1 = -5.468281666e-8
+ kt2 = -6.234897865e-02 lkt2 = 1.377966215e-8
+ at = 8.491634698e+04 lat = -2.313758535e-2
+ ute = -1.893419934e+00 lute = 8.446388674e-7
+ ua1 = -3.353153283e-09 lua1 = 2.920601073e-15 wua1 = 6.617444900e-30 pua1 = -3.308722450e-36
+ ub1 = 4.101751512e-18 lub1 = -3.204508915e-24 pub1 = 3.081487911e-45
+ uc1 = 3.188735465e-10 luc1 = -2.517695777e-16 wuc1 = -4.135903063e-31 puc1 = -2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.123 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.003044247e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.144612533e-9
+ k1 = 4.418300685e-01 lk1 = 3.390847368e-8
+ k2 = 1.155743619e-02 lk2 = -6.960452102e-09 wk2 = 1.387778781e-23 pk2 = -1.040834086e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.437694134e-01 ldsub = 2.314077213e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.743790865e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.671170052e-8
+ nfactor = {1.493771142e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.922958066e-7
+ eta0 = 4.153918492e-01 leta0 = 1.859720084e-8
+ etab = -1.234637215e-03 letab = 2.898534902e-10
+ u0 = 6.420346145e-03 lu0 = 1.070754753e-10
+ ua = -1.097309096e-09 lua = -5.157384327e-17
+ ub = 8.845879618e-19 lub = 1.755322802e-25
+ uc = -6.126448109e-11 luc = 1.502436844e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.347319152e+05 lvsat = -9.035390602e-3
+ a0 = 8.788192068e-01 la0 = -6.564572002e-8
+ ags = 9.950076829e-01 lags = 1.273087392e-7
+ a1 = 0.0
+ a2 = 1.106485264e+00 la2 = -7.738764019e-8
+ b0 = 1.751569461e-16 lb0 = -4.366049618e-23
+ b1 = 7.282076101e-20 lb1 = -1.815166699e-26
+ keta = -4.464049317e-02 lketa = 3.231132265e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.170588133e-01 lpclm = 2.877166222e-07 ppclm = -3.330669074e-28
+ pdiblc1 = -3.723560082e-01 lpdiblc1 = 1.936753674e-07 wpdiblc1 = 7.771561172e-22 ppdiblc1 = 1.387778781e-28
+ pdiblc2 = -8.352921763e-03 lpdiblc2 = 4.219915260e-09 wpdiblc2 = 5.204170428e-24 ppdiblc2 = 1.734723476e-30
+ pdiblcb = 2.163563710e-01 lpdiblcb = -1.257233392e-07 ppdiblcb = -1.110223025e-28
+ drout = 1.394365649e+00 ldrout = -2.157848363e-7
+ pscbe1 = 6.975643340e+08 lpscbe1 = 2.552696980e+1
+ pscbe2 = 2.047062388e-08 lpscbe2 = -2.897931263e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.545750116e+00 lbeta0 = 9.078136138e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.114932433e-12 lagidl = 5.566467413e-19
+ bgidl = 7.608364006e+08 lbgidl = 1.194060145e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.448437920e-01 lkt1 = 5.479659363e-9
+ kt2 = -1.673808726e-02 lkt2 = -8.992259540e-9
+ at = 9.344592137e+03 lat = 1.459274684e-2
+ ute = 4.294170626e-01 lute = -3.150723455e-7
+ ua1 = 4.691787198e-09 lua1 = -1.095956137e-15
+ ub1 = -4.457768141e-18 lub1 = 1.068959664e-24
+ uc1 = -2.726704746e-10 luc1 = 4.356764796e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.124 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.863580723e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.723039193e-8
+ k1 = -7.789825878e-01 lk1 = 3.382143405e-7
+ k2 = 5.505779462e-01 lk2 = -1.413193995e-07 wk2 = 2.220446049e-22 pk2 = 1.387778781e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.975951627e+00 ldsub = -2.969645439e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.269919322e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.202753912e-8
+ nfactor = {2.970405867e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.905988484e-7
+ eta0 = 1.128236100e+00 leta0 = -1.590899214e-7
+ etab = 6.456779281e-02 letab = -1.611238923e-08 wetab = -8.673617380e-25 petab = 7.155734338e-30
+ u0 = 1.161096607e-02 lu0 = -1.186764400e-9
+ ua = -5.772824102e-10 lua = -1.811982951e-16
+ ub = 1.690828730e-18 lub = -2.543532496e-26
+ uc = -1.080055805e-12 luc = 2.249767541e-20
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.561297911e+05 lvsat = -1.436913216e-2
+ a0 = -6.590336158e-01 la0 = 3.176871638e-7
+ ags = 2.160686824e+00 lags = -1.632542719e-7
+ a1 = 0.0
+ a2 = 1.161700591e+00 la2 = -9.115088873e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.120973870e-01 lketa = 2.004577490e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.761926159e-01 lpclm = -9.719195251e-9
+ pdiblc1 = 9.741129637e-01 lpdiblc1 = -1.419522208e-7
+ pdiblc2 = 2.117820294e-02 lpdiblc2 = -3.141160539e-9
+ pdiblcb = 9.751882474e-02 lpdiblcb = -9.610129823e-8
+ drout = -6.783329809e-01 ldrout = 3.008663877e-7
+ pscbe1 = 7.999049072e+08 lpscbe1 = 1.704682967e-2
+ pscbe2 = 1.304188057e-08 lpscbe2 = -1.046205562e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.033970329e+01 lbeta0 = -3.563883774e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.514075534e-12 lagidl = -9.867292966e-20
+ bgidl = 1.854155600e+09 lbgidl = -1.531201958e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.783538597e-01 lkt1 = -1.109395362e-8
+ kt2 = 4.941917831e-02 lkt2 = -2.548295034e-8
+ at = 1.406446700e+05 lat = -1.813576707e-2
+ ute = -2.757835876e+00 lute = 4.793982583e-7
+ ua1 = -7.754975894e-10 lua1 = 2.668466058e-16
+ ub1 = 5.361228676e-19 lub1 = -1.758425781e-25 pub1 = 3.851859889e-46
+ uc1 = -2.909190731e-10 luc1 = 4.811638486e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.125 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-8.131155341e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.513595908e-08 wvth0 = -1.734035738e-07 pvth0 = 3.403305242e-14
+ k1 = 3.790103419e-01 lk1 = 1.430142901e-07 wk1 = 6.166900660e-07 pk1 = -1.210346758e-13
+ k2 = -2.764987407e-01 lk2 = 7.605251241e-09 wk2 = 2.320907985e-09 pk2 = -4.555130057e-16
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.639517984e+00 ldsub = -4.553610397e-07 wdsub = -1.963558487e-06 pdsub = 3.853778065e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.229069174e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.778441566e-07 wvoff = 7.668797028e-07 pvoff = -1.505116449e-13
+ nfactor = {-2.418646791e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.179600709e-06 wnfactor = 5.086538381e-06 pnfactor = -9.983094554e-13
+ eta0 = 5.353696354e+00 leta0 = -1.003486642e-06 weta0 = -4.327122748e-06 peta0 = 8.492627461e-13
+ etab = 4.699172713e-01 letab = -9.719626947e-08 wetab = -4.191190945e-07 petab = 8.225840908e-14
+ u0 = -3.214105289e-02 lu0 = 7.287682747e-09 wu0 = 3.202691205e-08 pu0 = -6.285761894e-15
+ ua = -1.605103782e-08 lua = 2.838574974e-15 wua = 1.224018594e-14 pua = -2.402320094e-21
+ ub = 1.335519766e-17 lub = -2.317154768e-24 wub = -9.991776556e-24 pub = 1.961036026e-30
+ uc = -2.515553954e-10 luc = 4.918417369e-17 wuc = 2.120865029e-16 puc = -4.162515750e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.737661644e+05 lvsat = 4.901524870e-02 wvsat = 1.997880152e-01 pvsat = -3.921139480e-8
+ a0 = -3.728584921e+00 la0 = 9.502594562e-07 wa0 = 4.097602622e-06 pa0 = -8.042159787e-13
+ ags = 1.250000058e+00 lags = -9.593833283e-15
+ a1 = 0.0
+ a2 = 2.585973423e+00 la2 = -3.793297874e-07 wa2 = -1.635703518e-06 pa2 = 3.210313509e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.522196819e-01 lketa = 4.944785150e-08 wketa = 2.132236024e-07 pketa = -4.184833033e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.976049579e-01 lpclm = 4.783123892e-09 wpclm = 2.062519630e-08 ppclm = -4.048004152e-15
+ pdiblc1 = 3.681083740e+00 lpdiblc1 = -6.866974070e-07 wpdiblc1 = -2.961099865e-06 ppdiblc1 = 5.811602651e-13
+ pdiblc2 = -4.531180315e-02 lpdiblc2 = 9.610618995e-09 wpdiblc2 = 4.144182659e-08 ppdiblc2 = -8.133580095e-15
+ pdiblcb = -1.462075780e+01 lpdiblcb = 2.783467816e-06 wpdiblcb = 1.200255836e-05 ppdiblcb = -2.355682117e-12
+ drout = 1.000000945e+00 ldrout = -1.572365527e-13
+ pscbe1 = 8.000000007e+08 lpscbe1 = -1.211013794e-7
+ pscbe2 = -3.432331156e-08 lpscbe2 = 8.150710446e-15 wpscbe2 = 3.514658095e-14 ppscbe2 = -6.898043709e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.398125328e+00 lbeta0 = -9.121484305e-09 wbeta0 = -3.933440890e-08 pbeta0 = 7.719967762e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.817306669e-10 lagidl = -3.547823955e-17 wagidl = -1.529853045e-16 pagidl = 3.002566079e-23
+ bgidl = 1.000000285e+09 lbgidl = -4.730360031e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.493197995e+00 lkt1 = 1.870323723e-07 wkt1 = 8.065000661e-07 pkt1 = -1.582877355e-13
+ kt2 = 7.565266879e-01 lkt2 = -1.666799965e-07 wkt2 = -7.187388795e-07 pkt2 = 1.410632862e-13
+ at = -3.896816159e+05 lat = 8.422887629e-02 wat = 3.632023555e-01 pat = -7.128391031e-8
+ ute = -8.175028629e+00 lute = 1.588065733e-06 wute = 6.847879392e-06 pute = -1.343999049e-12
+ ua1 = -6.637865942e-09 lua1 = 1.442729841e-15 wua1 = 6.221177907e-15 pua1 = -1.220999482e-21
+ ub1 = 6.254904013e-18 lub1 = -1.314914606e-24 wub1 = -5.670028330e-24 pub1 = 1.112828110e-30
+ uc1 = -1.600035424e-10 luc1 = 2.698520553e-17 wuc1 = 1.163625807e-16 puc1 = -2.283790190e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.126 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.127 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.124648838e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.706194604e-7
+ k1 = 4.210818616e-01 lk1 = 2.114671972e-7
+ k2 = 2.113420949e-02 lk2 = 8.596014224e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = -1.694065895e-27 pcit = -1.761828530e-31
+ voff = {-2.804004741e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.598181832e-7
+ nfactor = {1.983803335e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.424216791e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.153077275e-02 lu0 = -2.044270362e-8
+ ua = -9.098047201e-10 lua = 1.854443048e-15
+ ub = 1.491779338e-18 lub = -5.043522411e-24
+ uc = -1.282516351e-10 luc = 4.517563002e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.672490943e+04 lvsat = 1.068582539e+0
+ a0 = 1.566615238e+00 la0 = -2.052229338e-6
+ ags = 6.394720045e-02 lags = 9.868197240e-7
+ a1 = 0.0
+ a2 = 1.083322921e+00 la2 = -2.266375124e-06 wa2 = -3.552713679e-21
+ b0 = -2.161420565e-07 lb0 = 1.728977587e-12
+ b1 = 9.955134135e-10 lb1 = -7.963375606e-15
+ keta = 4.018068624e-02 lketa = -3.363761825e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.896493835e-02 lpclm = 1.679237053e-06 wpclm = -5.551115123e-23 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.915673984e-03 lpdiblc2 = -1.276983438e-8
+ pdiblcb = -2.715826998e-01 lpdiblcb = 9.316197581e-7
+ drout = 0.56
+ pscbe1 = 8.000324970e+08 lpscbe1 = -6.499163959e-1
+ pscbe2 = 1.315044923e-08 lpscbe2 = -6.179421357e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.666054167e-11 lalpha0 = 1.333161838e-15
+ alpha1 = -6.666054167e-11 lalpha1 = 1.333161838e-15
+ beta0 = 4.581282086e+01 lbeta0 = -3.162447948e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.870274718e-09 lagidl = -1.939963340e-14 wagidl = 6.617444900e-30
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.235849912e-01 legidl = 1.047131499e-5
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365691544e-01 lkt1 = -3.361567574e-8
+ kt2 = -6.267063968e-02 lkt2 = 8.248976200e-8
+ at = 1.183123185e+05 lat = -9.464115887e-1
+ ute = -5.012560544e-02 lute = -6.570637432e-7
+ ua1 = 2.268500750e-09 lua1 = -3.565883958e-15
+ ub1 = -1.570875991e-18 lub1 = 6.839268476e-24
+ uc1 = -4.380619758e-11 luc1 = 2.803336491e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.128 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.069866256e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.239906809e-8
+ k1 = 4.556237202e-01 lk1 = -6.484228401e-8
+ k2 = 2.007683582e-02 lk2 = 1.705422642e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.164179846e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.199470589e-8
+ nfactor = {2.378038919e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.167837078e-06 wnfactor = -7.105427358e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.443397737e-03 lu0 = 4.254027232e-9
+ ua = -7.572954228e-10 lua = 6.344807637e-16
+ ub = 8.922232633e-19 lub = -2.475144842e-25 wub = -3.081487911e-39
+ uc = -7.084368051e-11 luc = -7.465141979e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.671623623e+05 lvsat = -8.547403617e-1
+ a0 = 1.370094967e+00 la0 = -4.802116133e-7
+ ags = 1.321801322e-01 lags = 4.410064215e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.426888399e-04 lketa = -8.219334060e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.401119263e-01 lpclm = -7.931506930e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.387319811e-03 lpdiblc2 = 1.365168829e-8
+ pdiblcb = -2.488330300e-01 lpdiblcb = 7.496391204e-7
+ drout = 0.56
+ pscbe1 = 1.224636900e+09 lpscbe1 = -3.397173053e+3
+ pscbe2 = -1.698011262e-08 lpscbe2 = 1.792281353e-13 ppscbe2 = 2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.446751046e+00 lbeta0 = 2.265262463e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.904539975e-10 lagidl = -1.962669803e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.670754974e+00 legidl = -6.281865390e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.063193317e-01 lkt1 = -2.755920237e-7
+ kt2 = -4.841666844e-02 lkt2 = -3.153153126e-8
+ at = -9.065933828e+04 lat = 7.252080717e-1
+ ute = -1.645263111e-01 lute = 2.580578176e-7
+ ua1 = 5.778773827e-10 lua1 = 9.957860376e-15
+ ub1 = 8.146409535e-19 lub1 = -1.224311373e-23
+ uc1 = -1.163111597e-11 luc1 = 2.295664482e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.129 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.063199473e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.736836213e-9
+ k1 = 4.427665361e-01 lk1 = -1.342299740e-8
+ k2 = 2.238297990e-02 lk2 = 7.831345119e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.585912374e-01 ldsub = -1.194145485e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.482687602e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.538498620e-8
+ nfactor = {9.059919706e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.719268760e-6
+ eta0 = 1.594707837e-01 leta0 = -3.178247240e-7
+ etab = -1.394757071e-01 letab = 2.778517638e-7
+ u0 = 8.601632881e-03 lu0 = 3.621202956e-9
+ ua = -7.352853466e-10 lua = 5.464566366e-16
+ ub = 8.528601283e-19 lub = -9.009087610e-26
+ uc = -7.556913799e-11 luc = 1.143321474e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.264314745e+00 la0 = -5.716847236e-8
+ ags = 1.560797535e-01 lags = 3.454255025e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.464757958e-03 lketa = -3.744375028e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.488073345e-01 lpclm = 2.361946495e-06 ppclm = 3.108624469e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.621872386e-03 lpdiblc2 = -6.381398745e-9
+ pdiblcb = -9.776424111e-02 lpdiblcb = 1.454750005e-7
+ drout = 0.56
+ pscbe1 = -4.171210305e+07 lpscbe1 = 1.667292191e+3
+ pscbe2 = 4.631193739e-08 lpscbe2 = -7.389354511e-14 ppscbe2 = 2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.144527102e+01 lbeta0 = -9.335576356e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.690680066e-10 lagidl = -2.774355581e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.815376811e-01 lkt1 = 2.522608815e-8
+ kt2 = -6.023855242e-02 lkt2 = 1.574731557e-8
+ at = 1.021557796e+05 lat = -4.591068088e-2
+ ute = -1.323451088e-01 lute = 1.293566616e-7
+ ua1 = 3.320607059e-09 lua1 = -1.011042424e-15
+ ub1 = -2.835183653e-18 lub1 = 2.353502076e-24
+ uc1 = 1.789645493e-11 luc1 = -9.513193603e-17 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.130 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.080253346e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.983204748e-8
+ k1 = 3.559763493e-01 lk1 = 1.600935854e-7
+ k2 = 5.664373486e-02 lk2 = -6.066498314e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.538016126e-01 ldsub = 1.029822606e-06 pdsub = -1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.107617634e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.985602103e-10
+ nfactor = {2.269123695e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.992787282e-9
+ eta0 = -2.188386675e-01 leta0 = 4.385161211e-07 weta0 = -2.151057110e-22 peta0 = -4.371503159e-28
+ etab = 8.242798594e-01 letab = -1.648951009e-06 wetab = 2.116362641e-22 petab = -9.436895709e-28
+ u0 = 1.231769894e-02 lu0 = -3.808197859e-9
+ ua = -2.809317911e-10 lua = -3.619165246e-16
+ ub = 9.337272840e-19 lub = -2.517657501e-25 wub = 3.081487911e-39
+ uc = -7.496753916e-11 luc = 1.023045924e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.949154737e+04 lvsat = -1.210264538e-2
+ a0 = 1.349266482e+00 la0 = -2.270095072e-7
+ ags = 1.615750419e-01 lags = 3.344389646e-7
+ a1 = 0.0
+ a2 = 6.001569927e-01 la2 = 3.995391301e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.083405178e-02 lketa = -2.858845418e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.592302506e-01 lpclm = 3.466122321e-7
+ pdiblc1 = 7.407420150e-01 lpdiblc1 = -7.012262346e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 1.203234000e-01 ldrout = 8.790300377e-7
+ pscbe1 = 7.981743154e+08 lpscbe1 = -1.186332945e+1
+ pscbe2 = 9.526279703e-09 lpscbe2 = -3.492672025e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.883960260e+00 lbeta0 = 1.782957602e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.471808281e-10 lagidl = 7.546826683e-16 pagidl = -8.271806126e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.587827164e-01 lkt1 = -2.026711633e-8
+ kt2 = -5.616202393e-02 lkt2 = 7.597254838e-9
+ at = 9.660944576e+04 lat = -3.482208970e-2
+ ute = 9.121531202e-01 lute = -1.958872090e-06 wute = 8.881784197e-22
+ ua1 = 6.057818692e-09 lua1 = -6.483453838e-15
+ ub1 = -4.209009179e-18 lub1 = 5.100143366e-24
+ uc1 = -1.262217768e-10 luc1 = 1.929986004e-16 wuc1 = -2.067951531e-31 puc1 = -2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.131 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.061395626e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.098818878e-8
+ k1 = 5.226190584e-01 lk1 = -6.426641356e-9
+ k2 = -5.745305410e-03 lk2 = 1.678201184e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.233157705e+00 ldsub = -4.560437967e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.128704363e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.505683220e-9
+ nfactor = {2.446759293e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.834978225e-7
+ eta0 = -1.229902487e-02 leta0 = 2.321282851e-7
+ etab = -1.649900875e+00 letab = 8.234112028e-7
+ u0 = 1.037583596e-02 lu0 = -1.867762149e-9
+ ua = -8.643992354e-11 lua = -5.562654406e-16
+ ub = 1.281983108e-19 lub = 5.531711593e-25
+ uc = -9.823827214e-11 luc = 3.348408823e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.177272666e+04 lvsat = 6.910189940e-02 pvsat = -1.164153218e-22
+ a0 = 1.496294625e+00 la0 = -3.739295848e-7
+ ags = -2.563720021e-01 lags = 7.520788176e-7
+ a1 = 0.0
+ a2 = 1.048426564e+00 la2 = -4.840096337e-8
+ b0 = -8.757847307e-17 lb0 = 8.751410289e-23
+ b1 = -3.641038050e-20 lb1 = 3.638361887e-26
+ keta = 1.074273877e-02 lketa = -2.441977703e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.551875389e+00 lpclm = -7.452298123e-7
+ pdiblc1 = 6.240057999e-02 lpdiblc1 = -2.338338057e-8
+ pdiblc2 = 7.601803479e-04 lpdiblc2 = -3.299376654e-10
+ pdiblcb = -1.455489873e-02 lpdiblcb = -1.043742412e-8
+ drout = 1.037783741e+00 ldrout = -3.775597026e-08 wdrout = -3.552713679e-21
+ pscbe1 = 8.238558016e+08 lpscbe1 = -3.752593977e+1
+ pscbe2 = 3.695351837e-09 lpscbe2 = 5.477374932e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.610435717e+00 lbeta0 = 1.057016105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.015367036e-09 lagidl = -5.069372234e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.243417019e-01 lkt1 = -5.468281666e-8
+ kt2 = -6.234897865e-02 lkt2 = 1.377966215e-8
+ at = 8.491634698e+04 lat = -2.313758535e-2
+ ute = -1.893419934e+00 lute = 8.446388674e-7
+ ua1 = -3.353153283e-09 lua1 = 2.920601073e-15 wua1 = 1.654361225e-30 pua1 = -1.654361225e-36
+ ub1 = 4.101751512e-18 lub1 = -3.204508915e-24 wub1 = -6.162975822e-39
+ uc1 = 3.188735465e-10 luc1 = -2.517695777e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.132 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.003044247e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.144612533e-9
+ k1 = 4.418300685e-01 lk1 = 3.390847368e-8
+ k2 = 1.155743619e-02 lk2 = -6.960452102e-09 wk2 = 1.387778781e-23 pk2 = 6.938893904e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.437694134e-01 ldsub = 2.314077213e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.743790865e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.671170052e-8
+ nfactor = {1.493771142e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.922958066e-7
+ eta0 = 4.153918492e-01 leta0 = 1.859720084e-8
+ etab = -1.234637215e-03 letab = 2.898534902e-10
+ u0 = 6.420346145e-03 lu0 = 1.070754753e-10
+ ua = -1.097309096e-09 lua = -5.157384327e-17
+ ub = 8.845879618e-19 lub = 1.755322802e-25
+ uc = -6.126448109e-11 luc = 1.502436844e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.347319152e+05 lvsat = -9.035390602e-3
+ a0 = 8.788192068e-01 la0 = -6.564572002e-8
+ ags = 9.950076829e-01 lags = 1.273087392e-7
+ a1 = 0.0
+ a2 = 1.106485264e+00 la2 = -7.738764019e-8
+ b0 = 1.751569461e-16 lb0 = -4.366049618e-23
+ b1 = 7.282076101e-20 lb1 = -1.815166699e-26
+ keta = -4.464049317e-02 lketa = 3.231132265e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.170588133e-01 lpclm = 2.877166222e-07 wpclm = 6.661338148e-22 ppclm = 1.110223025e-28
+ pdiblc1 = -3.723560082e-01 lpdiblc1 = 1.936753674e-07 wpdiblc1 = -1.665334537e-22 ppdiblc1 = -1.387778781e-29
+ pdiblc2 = -8.352921763e-03 lpdiblc2 = 4.219915260e-09 wpdiblc2 = 9.540979118e-24 ppdiblc2 = -2.818925648e-30
+ pdiblcb = 2.163563710e-01 lpdiblcb = -1.257233392e-07 wpdiblcb = 2.220446049e-22 ppdiblcb = 5.551115123e-29
+ drout = 1.394365649e+00 ldrout = -2.157848363e-7
+ pscbe1 = 6.975643340e+08 lpscbe1 = 2.552696980e+1
+ pscbe2 = 2.047062388e-08 lpscbe2 = -2.897931263e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.545750116e+00 lbeta0 = 9.078136138e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.114932433e-12 lagidl = 5.566467413e-19
+ bgidl = 7.608364006e+08 lbgidl = 1.194060145e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.448437920e-01 lkt1 = 5.479659363e-9
+ kt2 = -1.673808726e-02 lkt2 = -8.992259540e-9
+ at = 9.344592137e+03 lat = 1.459274684e-2
+ ute = 4.294170626e-01 lute = -3.150723455e-07 pute = 2.220446049e-28
+ ua1 = 4.691787198e-09 lua1 = -1.095956137e-15
+ ub1 = -4.457768141e-18 lub1 = 1.068959664e-24
+ uc1 = -2.726704746e-10 luc1 = 4.356764796e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.133 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.863580723e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.723039193e-8
+ k1 = -7.789825878e-01 lk1 = 3.382143405e-7
+ k2 = 5.505779462e-01 lk2 = -1.413193995e-07 wk2 = 8.881784197e-22 pk2 = 1.665334537e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.975951627e+00 ldsub = -2.969645439e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.269919322e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.202753912e-8
+ nfactor = {2.970405867e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.905988484e-7
+ eta0 = 1.128236100e+00 leta0 = -1.590899214e-7
+ etab = 6.456779281e-02 letab = -1.611238923e-08 wetab = 1.301042607e-23 petab = -1.214306433e-29
+ u0 = 1.161096607e-02 lu0 = -1.186764400e-9
+ ua = -5.772824102e-10 lua = -1.811982951e-16
+ ub = 1.690828730e-18 lub = -2.543532496e-26
+ uc = -1.080055805e-12 luc = 2.249767541e-20
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.561297911e+05 lvsat = -1.436913216e-2
+ a0 = -6.590336158e-01 la0 = 3.176871638e-7
+ ags = 2.160686824e+00 lags = -1.632542719e-7
+ a1 = 0.0
+ a2 = 1.161700591e+00 la2 = -9.115088873e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.120973870e-01 lketa = 2.004577490e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.761926159e-01 lpclm = -9.719195251e-9
+ pdiblc1 = 9.741129637e-01 lpdiblc1 = -1.419522208e-7
+ pdiblc2 = 2.117820294e-02 lpdiblc2 = -3.141160539e-9
+ pdiblcb = 9.751882474e-02 lpdiblcb = -9.610129823e-8
+ drout = -6.783329809e-01 ldrout = 3.008663877e-7
+ pscbe1 = 7.999049072e+08 lpscbe1 = 1.704682967e-2
+ pscbe2 = 1.304188057e-08 lpscbe2 = -1.046205562e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.033970329e+01 lbeta0 = -3.563883774e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.514075534e-12 lagidl = -9.867292966e-20
+ bgidl = 1.854155600e+09 lbgidl = -1.531201958e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.783538597e-01 lkt1 = -1.109395362e-8
+ kt2 = 4.941917831e-02 lkt2 = -2.548295034e-8
+ at = 1.406446700e+05 lat = -1.813576707e-2
+ ute = -2.757835876e+00 lute = 4.793982583e-7
+ ua1 = -7.754975894e-10 lua1 = 2.668466058e-16 pua1 = -4.135903063e-37
+ ub1 = 5.361228676e-19 lub1 = -1.758425781e-25 pub1 = -1.925929944e-46
+ uc1 = -2.909190731e-10 luc1 = 4.811638486e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.134 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-6.740392014e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.243177552e-08 wvth0 = -2.869332531e-07 pvth0 = 5.631495492e-14
+ k1 = 3.751617864e-01 lk1 = 1.437696268e-07 wk1 = 6.198316880e-07 pk1 = -1.216512662e-13
+ k2 = -4.549226187e-02 lk2 = -3.773323534e-08 wk2 = -1.862524528e-07 pk2 = 3.655483765e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.651771892e+00 ldsub = -4.577660530e-07 wdsub = -1.973561500e-06 pdsub = 3.873410477e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.229069217e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.778441650e-07 wvoff = 7.668797377e-07 pvoff = -1.505116517e-13
+ nfactor = {-2.418648291e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.179601003e-06 wnfactor = 5.086539606e-06 pnfactor = -9.983096957e-13
+ eta0 = 5.353695481e+00 leta0 = -1.003486470e-06 weta0 = -4.327122035e-06 peta0 = 8.492626062e-13
+ etab = 4.725328528e-01 letab = -9.770961656e-08 wetab = -4.212542250e-07 petab = 8.267746046e-14
+ u0 = -2.998961157e-02 lu0 = 6.865430115e-09 wu0 = 3.027066468e-08 pu0 = -5.941072004e-15
+ ua = -1.605103357e-08 lua = 2.838574139e-15 wua = 1.224018247e-14 pua = -2.402319413e-21
+ ub = 1.335527615e-17 lub = -2.317170172e-24 wub = -9.991840624e-24 pub = 1.961048600e-30
+ uc = -2.528789560e-10 luc = 4.944394231e-17 wuc = 2.131669413e-16 puc = -4.183720974e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.473416504e+05 lvsat = 4.382904146e-02 wvsat = 1.782173673e-01 pvsat = -3.497783159e-8
+ a0 = -3.728584082e+00 la0 = 9.502592916e-07 wa0 = 4.097601938e-06 pa0 = -8.042158443e-13
+ ags = 1.250000058e+00 lags = -9.593840389e-15
+ a1 = 0.0
+ a2 = 2.596181299e+00 la2 = -3.813332362e-07 wa2 = -1.644036329e-06 pa2 = 3.226667902e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.522196895e-01 lketa = 4.944785299e-08 wketa = 2.132236087e-07 pketa = -4.184833155e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.974762430e-01 lpclm = 4.808386125e-09 wpclm = 2.073026783e-08 ppclm = -4.068626016e-15
+ pdiblc1 = 3.699562970e+00 lpdiblc1 = -6.903242329e-07 wpdiblc1 = -2.976184682e-06 ppdiblc1 = 5.841208866e-13
+ pdiblc2 = -4.557042767e-02 lpdiblc2 = 9.661377936e-09 wpdiblc2 = 4.165294488e-08 ppdiblc2 = -8.175015227e-15
+ pdiblcb = -1.469566173e+01 lpdiblcb = 2.798168836e-06 wpdiblcb = 1.206370334e-05 ppdiblcb = -2.367682737e-12
+ drout = 1.000000945e+00 ldrout = -1.572365740e-13 wdrout = -8.526512829e-20 pdrout = 1.776356839e-26
+ pscbe1 = 8.000000007e+08 lpscbe1 = -1.211013794e-7
+ pscbe2 = -3.454264956e-08 lpscbe2 = 8.193758818e-15 wpscbe2 = 3.532562919e-14 ppscbe2 = -6.933184613e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.398370801e+00 lbeta0 = -9.169662029e-09 wbeta0 = -3.953479131e-08 pbeta0 = 7.759295817e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.022247156e-10 lagidl = -1.987400402e-17 wagidl = -8.808364242e-17 pagidl = 1.728773608e-23
+ bgidl = 1.000000285e+09 lbgidl = -4.730360031e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.493197741e+00 lkt1 = 1.870323226e-07 wkt1 = 8.064998591e-07 pkt1 = -1.582876948e-13
+ kt2 = 7.610120957e-01 lkt2 = -1.675603251e-07 wkt2 = -7.224003718e-07 pkt2 = 1.417819090e-13
+ at = -3.919482398e+05 lat = 8.467373522e-02 wat = 3.650526278e-01 pat = -7.164705399e-8
+ ute = -8.217763943e+00 lute = 1.596453180e-06 wute = 6.882764742e-06 pute = -1.350845822e-12
+ ua1 = -6.676690223e-09 lua1 = 1.450349688e-15 wua1 = 6.252870633e-15 pua1 = -1.227219655e-21
+ ub1 = 6.290288754e-18 lub1 = -1.321859392e-24 wub1 = -5.698913319e-24 pub1 = 1.118497223e-30
+ uc1 = -1.607297221e-10 luc1 = 2.712772920e-17 wuc1 = 1.169553700e-16 puc1 = -2.295424568e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.135 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.136 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.185320336e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.684004831e-06 wvth0 = 4.710001210e-08 pvth0 = -9.419656235e-13
+ k1 = 4.791227057e-01 lk1 = -9.493070259e-07 wk1 = -4.505780381e-08 pk1 = 9.011229587e-13
+ k2 = -2.750372412e-02 lk2 = 9.813189376e-07 wk2 = 3.775821152e-08 pk2 = -7.551364781e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = -3.388131789e-27 pcit = 3.388131789e-32
+ voff = {-4.477709590e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.807104865e-06 wvoff = 1.299317159e-07 pvoff = -2.598538818e-12
+ nfactor = {-9.118769647e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.789723549e-05 wnfactor = 2.247951364e-06 pnfactor = -4.495737505e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.725450538e-02 lu0 = -1.349131495e-07 wu0 = -4.443402332e-09 pu0 = 8.886478075e-14
+ ua = -7.382989945e-10 lua = -1.575545406e-15 wua = -1.331419528e-16 pua = 2.662741196e-21
+ ub = 1.073058464e-18 lub = 3.330587315e-24 wub = 3.250580393e-25 pub = -6.500921869e-30
+ uc = -4.709998077e-10 luc = 7.306467832e-15 wuc = 2.660795194e-16 puc = -5.321394819e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.343008928e+05 lvsat = 2.028839223e+01 wvsat = 7.460558626e-01 pvsat = -1.492056890e-5
+ a0 = 7.034262548e-01 la0 = 1.521091588e-05 wa0 = 6.701039659e-07 pa0 = -1.340158679e-11
+ ags = -6.449066257e-01 lags = 1.516337524e-05 wags = 5.502917315e-07 pags = -1.100543017e-11
+ a1 = 0.0
+ a2 = 1.083322921e+00 la2 = -2.266375124e-6
+ b0 = 5.803974115e-08 lb0 = -3.754456842e-12 wb0 = -2.128506197e-13 pb0 = 4.256855948e-18
+ b1 = 9.346462525e-09 lb1 = -1.749762199e-13 wb1 = -6.482942007e-15 pb1 = 1.296540752e-19
+ keta = 1.273353118e-01 lketa = -2.079404635e-06 wketa = -6.765918167e-08 pketa = 1.353133904e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.896493835e-02 lpclm = 1.679237053e-06 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.031147370e-03 lpdiblc2 = -1.507921721e-08 wpdiblc2 = -8.964337467e-11 ppdiblc2 = 1.792801606e-15
+ pdiblcb = -9.482541773e-01 lpdiblcb = 1.446455195e-05 wpdiblcb = 5.253081880e-07 ppdiblcb = -1.050577766e-11
+ drout = 0.56
+ pscbe1 = 8.005045564e+08 lpscbe1 = -1.009075794e+01 wpscbe1 = -3.664653968e-01 ppscbe1 = 7.329038583e-6
+ pscbe2 = 7.541066414e-08 lpscbe2 = -1.306952751e-12 wpscbe2 = -4.833335196e-14 ppscbe2 = 9.666315142e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.666054167e-11 lalpha0 = 1.333161838e-15
+ alpha1 = -6.666054167e-11 lalpha1 = 1.333161838e-15
+ beta0 = 1.406535457e+01 lbeta0 = 3.186811965e-04 wbeta0 = 2.464593905e-05 pbeta0 = -4.929006662e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.757549771e-09 lagidl = -3.714448231e-14 wagidl = -6.888022708e-16 pagidl = 1.377553915e-20
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -8.029306234e+00 legidl = 1.625801496e-04 wegidl = 5.904412669e-06 pegidl = -1.180839136e-10
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.232094334e-01 lkt1 = -2.300726777e-06 wkt1 = -8.800251176e-08 pkt1 = 1.759985553e-12
+ kt2 = -2.588107810e-02 lkt2 = -6.532744293e-07 wkt2 = -2.856017813e-08 pkt2 = 5.711825708e-13
+ at = 7.163679682e+05 lat = -1.290708501e+01 wat = -4.642777775e-01 pat = 9.285214306e-6
+ ute = -8.918971645e+00 lute = 1.767133385e-04 wute = 6.884991607e-06 pute = -1.376947717e-10
+ ua1 = -1.954914943e-08 lua1 = 4.327710837e-13 wua1 = 1.693730365e-14 pua1 = -3.387336240e-19
+ ub1 = 1.402668815e-17 lub1 = -3.051005502e-22 wub1 = -1.210857622e-23 pub1 = 2.421626245e-28
+ uc1 = 6.890242163e-10 luc1 = -1.437573600e-14 wuc1 = -5.689050442e-16 puc1 = 1.137768274e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.137 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.962411700e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.715104755e-07 wvth0 = -5.715603750e-08 pvth0 = -1.079938549e-13
+ k1 = 3.866964278e-01 lk1 = -2.099647355e-07 wk1 = 5.350908429e-08 pk1 = 1.126603006e-13
+ k2 = 7.010276894e-02 lk2 = 2.005387339e-07 wk2 = -3.883573219e-08 pk2 = -1.424412250e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {3.103787478e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.257535550e-06 wvoff = -4.089586249e-07 pvoff = 1.712187824e-12
+ nfactor = {2.118417299e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.188549236e-04 wnfactor = -1.459942755e-05 pnfactor = 8.980927348e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.554659554e-03 lu0 = -7.332004219e-08 wu0 = -8.626858836e-10 pu0 = 6.022168098e-14
+ ua = 1.015514733e-09 lua = -1.560476617e-14 wua = -1.376253798e-15 pua = 1.260672227e-20
+ ub = 3.317841857e-19 lub = 9.260236706e-24 wub = 4.350755813e-25 pub = -7.380981342e-30
+ uc = 4.544893604e-10 luc = -9.676527836e-17 wuc = -4.078223436e-16 puc = 6.932476747e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.226675710e+06 lvsat = -1.299636227e+01 wvsat = -2.297505726e+00 pvsat = 9.425686791e-6
+ a0 = 4.283772827e+00 la0 = -1.342922514e-05 wa0 = -2.261923087e-06 pa0 = 1.005247459e-11
+ ags = 1.395879712e+00 lags = -1.161415487e-06 wags = -9.810251485e-07 pags = 1.243979357e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -2.766479371e-07 lb0 = -1.077201411e-12 wb0 = 2.147651134e-13 pb0 = 8.362443817e-19
+ b1 = -3.911180911e-08 lb1 = 2.126543363e-13 wb1 = 3.036296675e-14 pb1 = -1.650861132e-19
+ keta = -1.225815475e-01 lketa = -8.025344911e-08 wketa = 9.450733687e-08 pketa = 5.592094792e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.649027600e+00 lpclm = -7.605756053e-05 wpclm = -7.304254145e-06 ppclm = 5.842866453e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -2.491669213e-02 lpdiblc2 = 2.004836921e-07 wpdiblc2 = 1.826613408e-08 ppdiblc2 = -1.450399266e-13
+ pdiblcb = -5.950373434e-01 lpdiblcb = 1.163907690e-05 wpdiblcb = 2.687625630e-07 ppdiblcb = -8.453601219e-12
+ drout = 0.56
+ pscbe1 = 7.393014417e+09 lpscbe1 = -5.274532415e+04 wpscbe1 = -4.788585487e+03 ppscbe1 = 3.830956187e-2
+ pscbe2 = -4.759839385e-07 lpscbe2 = 3.103798795e-12 wpscbe2 = 3.563301781e-13 ppscbe2 = -2.270379298e-18
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.352357080e-09 lalpha0 = 1.161778916e-14 walpha0 = 1.127482230e-15 palpha0 = -9.019029139e-21
+ alpha1 = -1.352357080e-09 lalpha1 = 1.161778916e-14 walpha1 = 1.127482230e-15 palpha1 = -9.019029139e-21
+ beta0 = 4.020727757e+02 lbeta0 = -2.785092987e-03 wbeta0 = -3.094581664e-04 pbeta0 = 2.179686611e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.435528843e-10 lagidl = -1.223479600e-14 wagidl = 3.640989696e-17 pagidl = 7.974374835e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 2.448791870e+01 legidl = -9.753374969e-05 wegidl = -1.771323801e-05 pegidl = 7.083993280e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.964582714e-01 lkt1 = -2.514716411e-06 wkt1 = -8.528645950e-08 pkt1 = 1.738259132e-12
+ kt2 = -1.913907696e-01 lkt2 = 6.706814534e-07 wkt2 = 1.109925104e-07 pkt2 = -5.451363665e-13
+ at = -1.735030178e+06 lat = 6.702298381e+00 wat = 1.276544815e+00 pat = -4.640086932e-6
+ ute = 2.523684590e+01 lute = -9.650809741e-05 wute = -1.971939007e-05 pute = 7.512072750e-11
+ ua1 = 5.183258511e-08 lua1 = -1.382303270e-13 wua1 = -3.978964466e-14 pua1 = 1.150402681e-19
+ ub1 = -2.974360404e-17 lub1 = 4.502961616e-23 wub1 = 2.372273229e-23 pub1 = -4.446150749e-29
+ uc1 = -8.197451350e-09 luc1 = 5.670953697e-14 wuc1 = 6.354750478e-15 puc1 = -4.400647255e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.138 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.156853555e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.506535739e-07 wvth0 = -1.145169793e-07 pvth0 = 1.214077520e-13
+ k1 = 1.266264686e+00 lk1 = -3.727591286e-06 wk1 = -6.392914959e-07 pk1 = 2.883353413e-12
+ k2 = -2.138588179e-01 lk2 = 1.336176369e-06 wk2 = 1.833973425e-07 pk2 = -1.031210182e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.397288766e-01 ldsub = -1.118709906e-06 wdsub = 1.464307701e-08 pdsub = -5.856154539e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-4.484586270e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.772562035e-07 wvoff = 1.554097959e-07 pvoff = -5.448710484e-13
+ nfactor = {-1.936693999e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.331972331e-05 wnfactor = 1.573812036e-05 pnfactor = -3.151862007e-11
+ eta0 = 1.594707837e-01 leta0 = -3.178247240e-7
+ etab = -1.394938409e-01 letab = 2.779242858e-07 wetab = 1.407752314e-11 petab = -5.629974557e-17
+ u0 = -4.059792307e-02 lu0 = 1.272534262e-07 wu0 = 3.819420568e-08 pu0 = -9.597717847e-14
+ ua = -9.500179521e-09 lua = 2.645028181e-14 wua = 6.804292526e-15 pua = -2.010945033e-20
+ ub = 5.266294080e-18 lub = -1.047417601e-23 wub = -3.426201738e-24 pub = 8.061289896e-30
+ uc = 7.658259362e-10 luc = -1.341882749e-15 wuc = -6.531850929e-16 puc = 1.050595423e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -3.845227433e+05 lvsat = 1.445777308e+00 wvsat = 3.399941805e-01 pvsat = -1.122374273e-6
+ a0 = -6.954349099e-01 la0 = 6.483946087e-06 wa0 = 1.521377174e-06 pa0 = -5.077945726e-12
+ ags = 3.027560770e+00 lags = -7.686940434e-06 wags = -2.229165171e-06 pags = 6.235622065e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -2.642922917e-07 lb0 = -1.126614911e-12 wb0 = 2.051732776e-13 pb0 = 8.746046749e-19
+ b1 = 3.740708951e-08 lb1 = -9.336501675e-14 wb1 = -2.903957247e-14 pb1 = 7.248038288e-20
+ keta = -2.281824881e-01 lketa = 3.420726965e-07 wketa = 1.821594729e-07 pketa = -2.946231718e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.733823673e+01 lpclm = 3.187166117e-05 wpclm = 1.303383552e-05 ppclm = -2.290874562e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 5.015220661e-02 lpdiblc2 = -9.973672719e-08 wpdiblc2 = -3.612205682e-08 ppdiblc2 = 7.247286173e-14
+ pdiblcb = 4.654673250e+00 lpdiblcb = -9.355906941e-06 wpdiblcb = -3.689374254e-06 ppdiblcb = 7.376036818e-12
+ drout = 0.56
+ pscbe1 = -1.226862412e+10 lpscbe1 = 2.588677871e+04 wpscbe1 = 9.491898524e+03 ppscbe1 = -1.880187802e-2
+ pscbe2 = 5.924246864e-07 lpscbe2 = -1.169050424e-12 wpscbe2 = -4.239538804e-13 ppscbe2 = 8.501834267e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.004714161e-09 lalpha0 = -5.807293356e-15 walpha0 = -2.254964460e-15 palpha0 = 4.508271520e-21
+ alpha1 = 3.004714161e-09 lalpha1 = -5.807293356e-15 walpha1 = -2.254964460e-15 palpha1 = 4.508271520e-21
+ beta0 = -6.128613637e+02 lbeta0 = 1.273897594e-03 wbeta0 = 4.846567322e-04 pbeta0 = -9.961893090e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 5.166263542e-09 lagidl = -3.032231444e-14 wagidl = -3.801751660e-15 pagidl = 2.332420002e-20
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.148357657e+00 lkt1 = 8.922549863e-07 wkt1 = 5.176603494e-07 pkt1 = -6.730849380e-13
+ kt2 = -1.786909774e-02 lkt2 = -2.327769579e-08 wkt2 = -3.289191610e-08 pkt2 = 3.029558462e-14
+ at = -7.659297368e+05 lat = 2.826608905e+00 wat = 6.739052034e-01 pat = -2.229971425e-6
+ ute = -7.090644051e-01 lute = 7.256473579e-06 wute = 4.477141103e-07 pute = -5.532866389e-12
+ ua1 = 9.758585284e-09 lua1 = 3.003474786e-14 wua1 = -4.997879752e-15 pua1 = -2.410121955e-20
+ ub1 = -1.648499006e-17 lub1 = -7.995094686e-24 wub1 = 1.059650851e-23 pub1 = 8.033739849e-30
+ uc1 = 1.293950600e-08 luc1 = -2.782275675e-14 wuc1 = -1.003120055e-14 puc1 = 2.152528787e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.139 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.963605242e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.063746725e-08 wvth0 = -6.512700396e-08 pvth0 = 2.266410297e-14
+ k1 = -1.830332532e+00 lk1 = 2.463327151e-06 wk1 = 1.697257821e-06 pk1 = -1.788027856e-12
+ k2 = 9.110662651e-01 lk2 = -9.128469765e-07 wk2 = -6.632984633e-07 pk2 = 6.615591077e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -7.717407440e+00 ldsub = 1.598927323e-05 wdsub = 5.794086767e-06 pdsub = -1.161320103e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.687384880e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.180215199e-07 wvoff = -3.262317291e-08 pvoff = -1.689433151e-13
+ nfactor = {2.650602277e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -6.991783369e-07 wnfactor = -2.961464006e-07 pnfactor = 5.381282604e-13
+ eta0 = 3.700363400e+00 leta0 = -7.397007401e-06 weta0 = -3.042523596e-06 peta0 = 6.082810936e-12
+ etab = 1.279438731e+01 letab = -2.558033161e-05 wetab = -9.292538053e-06 petab = 1.857821793e-11
+ u0 = 3.989827779e-02 lu0 = -3.367981085e-08 wu0 = -2.141113433e-08 pu0 = 2.318969163e-14
+ ua = 5.452434252e-09 lua = -3.443955567e-15 wua = -4.450880859e-15 pua = 2.392623893e-21
+ ub = 2.040095213e-18 lub = -4.024149529e-24 wub = -8.588866997e-25 pub = 2.928546796e-30
+ uc = 5.608126623e-10 luc = -9.320068863e-16 wuc = -4.935637998e-16 puc = 7.314701582e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.940097215e+05 lvsat = -7.104949004e-01 wvsat = -4.925840728e-01 pvsat = 5.421702883e-7
+ a0 = 5.933972780e+00 la0 = -6.769996677e-06 wa0 = -3.559162515e-06 pa0 = 5.079399456e-12
+ ags = -1.142733332e+00 lags = 6.505826048e-07 wags = 1.012550242e-06 pags = -2.454261016e-13
+ a1 = 0.0
+ a2 = -2.302810494e+00 la2 = 6.203340423e-06 wa2 = 2.253608496e-06 pa2 = -4.505560589e-12
+ b0 = -1.174249786e-06 lb0 = 6.926312589e-13 wb0 = 9.115841999e-13 pb0 = -5.376979578e-19
+ b1 = -6.965714733e-08 lb1 = 1.206847647e-13 wb1 = 5.407567936e-14 pb1 = -9.368903107e-20
+ keta = 8.330025912e-02 lketa = -2.806638581e-07 wketa = -7.307759516e-08 pketa = 2.156633650e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.182002613e+00 lpclm = 9.567392758e-06 wpclm = 5.155668767e-06 ppclm = -7.158202571e-12
+ pdiblc1 = 5.753534132e+00 lpdiblc1 = -1.072312607e-05 wpdiblc1 = -3.891490674e-06 ppdiblc1 = 7.780121102e-12
+ pdiblc2 = 1.011402042e-04 lpdiblc2 = 3.286180838e-10 wpdiblc2 = 2.552978058e-10 ppdiblc2 = -2.551101619e-16
+ pdiblcb = -2.928112643e+00 lpdiblcb = 5.804091498e-06 wpdiblcb = 2.253721182e-06 ppdiblcb = -4.505785879e-12
+ drout = -3.706480286e+00 ldrout = 8.529824708e-06 wdrout = 2.970793623e-06 pdrout = -5.939403712e-12
+ pscbe1 = 7.716539830e+08 lpscbe1 = -1.841929003e+02 wpscbe1 = 2.058805231e+01 ppscbe1 = 1.337815138e-4
+ pscbe2 = 6.097189690e-09 lpscbe2 = 3.173618998e-15 wpscbe2 = 2.662043726e-15 ppscbe2 = -2.734858832e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.358864408e+01 lbeta0 = 1.465369324e-06 wbeta0 = -1.374435850e-05 pbeta0 = 2.465475917e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -9.962258505e-09 lagidl = -7.638981238e-17 wagidl = 7.541931381e-15 pagidl = 6.451715396e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.249036580e-01 lkt1 = 4.455112264e-07 wkt1 = 3.618552804e-07 pkt1 = -3.615893168e-13
+ kt2 = -1.047926747e-02 lkt2 = -3.805192479e-08 wkt2 = -3.546407203e-08 pkt2 = 3.543800594e-14
+ at = 1.088440409e+06 lat = -8.807684255e-01 wat = -7.699702791e-01 pat = 6.567182918e-7
+ ute = 6.886255334e+00 lute = -7.928583339e-06 wute = -4.637767238e-06 pute = 4.634358479e-12
+ ua1 = 4.997483351e-08 lua1 = -5.036818965e-14 wua1 = -3.409330561e-14 pua1 = 3.406824703e-20
+ ub1 = -4.242780867e-17 lub1 = 4.387147457e-23 wub1 = 2.966971267e-23 pub1 = -3.009864967e-29
+ uc1 = -2.020124890e-09 luc1 = 2.085509695e-15 wuc1 = 1.470259713e-15 puc1 = -1.469179073e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.140 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.521224666e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.356807539e-08 wvth0 = -8.483006529e-08 pvth0 = 4.235268255e-14
+ k1 = 7.596823015e-01 lk1 = -1.247840214e-07 wk1 = -1.840350404e-07 pk1 = 9.188225444e-14
+ k2 = -2.520232930e-03 lk2 = 6.803537281e-11 wk2 = -2.503662467e-09 pk2 = 1.249991042e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.623581880e+01 ldsub = -7.946347390e-06 wdsub = -1.164674584e-05 pdsub = 5.814812563e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {3.063602595e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.567280301e-07 wvoff = -4.030850199e-07 pvoff = 2.012462425e-13
+ nfactor = {1.822784583e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.280309109e-07 wnfactor = 4.843990548e-07 pnfactor = -2.418434941e-13
+ eta0 = -7.850703160e+00 leta0 = 4.145569126e-06 weta0 = 6.085047191e-06 peta0 = -3.038051086e-12
+ etab = -2.559004323e+01 letab = 1.277588638e-05 wetab = 1.858501980e-05 petab = -9.278849908e-12
+ u0 = 5.753224219e-03 lu0 = 4.401461039e-10 wu0 = 3.588588969e-09 pu0 = -1.791656872e-15
+ ua = 5.207786029e-09 lua = -3.199487161e-15 wua = -4.109971138e-15 pua = 2.051964740e-21
+ ub = -5.205459750e-18 lub = 3.216079951e-24 wub = 4.140582757e-24 pub = -2.067248050e-30
+ uc = -7.120871571e-10 luc = 3.399573518e-16 wuc = 4.765382556e-16 puc = -2.379188722e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.504536300e+05 lvsat = 1.333477706e-01 wvsat = 9.989652945e-02 pvsat = -4.987484077e-8
+ a0 = -2.427006638e+00 la0 = 1.584837420e-06 wa0 = 3.045705850e-06 pa0 = -1.520614331e-12
+ ags = -2.230784136e+00 lags = 1.737833692e-06 wags = 1.532759833e-06 pags = -7.652533378e-13
+ a1 = 0.0
+ a2 = 6.854361538e+00 la2 = -2.947101088e-06 wa2 = -4.507216992e-06 pa2 = 2.250295691e-12
+ b0 = -9.615109074e-07 lb0 = 4.800487432e-13 wb0 = 7.464324554e-13 pb0 = -3.726675999e-19
+ b1 = 1.021576308e-07 lb1 = -5.100372953e-14 wb1 = -7.930619467e-14 pb1 = 3.959480728e-20
+ keta = -3.567370423e-01 lketa = 1.590500159e-07 wketa = 2.852789638e-07 pketa = -1.424298019e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.720733326e+00 lpclm = -3.325859670e-06 wpclm = -4.012646442e-06 ppclm = 2.003373926e-12
+ pdiblc1 = -9.963183654e+00 lpdiblc1 = 4.982039932e-06 wpdiblc1 = 7.782981348e-06 ppdiblc1 = -3.885770182e-12
+ pdiblc2 = 7.601803479e-04 lpdiblc2 = -3.299376654e-10
+ pdiblcb = 5.791670387e+00 lpdiblcb = -2.909282491e-06 wpdiblcb = -4.507442364e-06 ppdiblcb = 2.250408212e-12
+ drout = 8.691391112e+00 ldrout = -3.858934254e-06 wdrout = -5.941587245e-06 pdrout = 2.966426556e-12
+ pscbe1 = 4.261949799e+08 lpscbe1 = 1.610121904e+02 wpscbe1 = 3.087088678e+02 ppscbe1 = -1.541275329e-4
+ pscbe2 = 3.887984973e-09 lpscbe2 = 5.381199949e-15 wpscbe2 = -1.495434153e-16 ppscbe2 = 7.466179324e-23
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.135860091e+01 lbeta0 = -1.629152659e-05 wbeta0 = -2.697541761e-05 pbeta0 = 1.346788188e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.006265211e-08 lagidl = 1.001658001e-14 wagidl = 1.636311920e-14 pagidl = -8.169532709e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.243417019e-01 lkt1 = -5.468281666e-8
+ kt2 = -6.234897865e-02 lkt2 = 1.377966215e-8
+ at = 3.752276113e+05 lat = -1.680798387e-01 wat = -2.253721182e-01 pat = 1.125204106e-7
+ ute = -1.893419934e+00 lute = 8.446388674e-7
+ ua1 = -3.353153283e-09 lua1 = 2.920601073e-15 wua1 = -1.654361225e-30 pua1 = -2.481541838e-36
+ ub1 = 5.262996569e-18 lub1 = -3.784277929e-24 wub1 = -9.014884728e-25 pub1 = 4.500816424e-31
+ uc1 = 3.188735465e-10 luc1 = -2.517695777e-16 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.141 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.003044247e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.144612533e-9
+ k1 = 4.418300685e-01 lk1 = 3.390847368e-8
+ k2 = 1.155743619e-02 lk2 = -6.960452102e-09 wk2 = 1.387778781e-23 pk2 = 1.734723476e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.437694134e-01 ldsub = 2.314077213e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.743790865e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.671170052e-8
+ nfactor = {1.493771142e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.922958066e-7
+ eta0 = 4.153918492e-01 leta0 = 1.859720084e-8
+ etab = -1.234637215e-03 letab = 2.898534902e-10
+ u0 = 6.420346145e-03 lu0 = 1.070754753e-10
+ ua = -1.097309096e-09 lua = -5.157384327e-17
+ ub = 8.845879618e-19 lub = 1.755322802e-25
+ uc = -6.126448109e-11 luc = 1.502436844e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.347319152e+05 lvsat = -9.035390602e-3
+ a0 = 8.788192068e-01 la0 = -6.564572002e-8
+ ags = 9.950076829e-01 lags = 1.273087392e-7
+ a1 = 0.0
+ a2 = 1.106485264e+00 la2 = -7.738764019e-8
+ b0 = 1.751569461e-16 lb0 = -4.366049618e-23
+ b1 = 7.282076101e-20 lb1 = -1.815166699e-26
+ keta = -4.464049317e-02 lketa = 3.231132265e-09 wketa = 1.110223025e-22
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.170588133e-01 lpclm = 2.877166222e-07 wpclm = -2.220446049e-22 ppclm = -2.220446049e-28
+ pdiblc1 = -3.723560082e-01 lpdiblc1 = 1.936753674e-07 wpdiblc1 = 3.885780586e-22 ppdiblc1 = -1.249000903e-28
+ pdiblc2 = -8.352921763e-03 lpdiblc2 = 4.219915260e-09 wpdiblc2 = -4.770489559e-24 ppdiblc2 = -2.710505431e-30
+ pdiblcb = 2.163563710e-01 lpdiblcb = -1.257233392e-07 wpdiblcb = 1.110223025e-22 ppdiblcb = -5.551115123e-29
+ drout = 1.394365649e+00 ldrout = -2.157848363e-7
+ pscbe1 = 6.975643340e+08 lpscbe1 = 2.552696980e+1
+ pscbe2 = 2.047062388e-08 lpscbe2 = -2.897931263e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.545750116e+00 lbeta0 = 9.078136138e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.114932433e-12 lagidl = 5.566467413e-19
+ bgidl = 7.608364006e+08 lbgidl = 1.194060145e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.448437920e-01 lkt1 = 5.479659363e-9
+ kt2 = -1.673808726e-02 lkt2 = -8.992259540e-9
+ at = 9.344592137e+03 lat = 1.459274684e-2
+ ute = 4.294170626e-01 lute = -3.150723455e-7
+ ua1 = 4.691787198e-09 lua1 = -1.095956137e-15
+ ub1 = -4.457768141e-18 lub1 = 1.068959664e-24
+ uc1 = -2.726704746e-10 luc1 = 4.356764796e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.142 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-7.148446706e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.998268001e-08 wvth0 = -1.331479119e-07 pvth0 = 3.318911426e-14
+ k1 = -2.117888029e+00 lk1 = 6.719566052e-07 wk1 = 1.039408361e-06 pk1 = -2.590881250e-13
+ k2 = 1.560399840e+00 lk2 = -3.930326540e-07 wk2 = -7.839368543e-07 pk2 = 1.954080200e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.239072385e+00 ldsub = -1.359611340e-06 wdsub = -3.309511801e-06 pdsub = 8.249454592e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.675794140e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.575385228e-07 wvoff = 1.275554324e-06 pvoff = -3.179510487e-13
+ nfactor = {-1.060119757e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.307148183e-06 wnfactor = 8.460433062e-06 pnfactor = -2.108889847e-12
+ eta0 = 1.039940686e+01 leta0 = -2.470068301e-06 weta0 = -7.197321114e-06 peta0 = 1.794040248e-12
+ etab = 9.745245310e-01 letab = -2.429327556e-07 wetab = -7.064103353e-07 petab = 1.760833722e-13
+ u0 = -5.548715835e-02 lu0 = 1.553844958e-08 wu0 = 5.208907916e-08 pu0 = -1.298398432e-14
+ ua = -2.680275910e-08 lua = 6.355895153e-15 wua = 2.035915226e-14 pua = -5.074824089e-21
+ ub = 2.309902216e-17 lub = -5.361748660e-24 wub = -1.661943746e-23 pub = 4.142644078e-30
+ uc = -4.615441086e-10 luc = 1.148000698e-16 wuc = 3.574637697e-16 puc = -8.910320656e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.326580675e+05 lvsat = 5.761557344e-02 wvsat = 2.241894801e-01 pvsat = -5.588259077e-8
+ a0 = -9.438434903e+00 la0 = 2.506084626e-06 wa0 = 6.815554572e-06 pa0 = -1.698879210e-12
+ ags = 2.160686814e+00 lags = -1.632542695e-07 wags = 7.556565151e-15 pags = -1.883586620e-21
+ a1 = 0.0
+ a2 = 4.713000355e+00 la2 = -9.763656243e-07 wa2 = -2.756916622e-06 pa2 = 6.872028218e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.689450355e-01 lketa = 1.339219040e-07 wketa = 3.546563117e-07 pketa = -8.840340554e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.314135251e-01 lpclm = 1.442664801e-09 wpclm = 3.476254549e-08 ppclm = -8.665085901e-15
+ pdiblc1 = 7.403002208e+00 lpdiblc1 = -1.744449298e-06 wpdiblc1 = -4.990823867e-06 ppdiblc1 = 1.244037711e-12
+ pdiblc2 = -6.879670003e-02 lpdiblc2 = 1.928643365e-08 wpdiblc2 = 6.984859688e-08 ppdiblc2 = -1.741081050e-14
+ pdiblcb = -2.596140478e+01 lpdiblcb = 6.399476293e-06 wpdiblcb = 2.022985510e-05 ppdiblcb = -5.042594831e-12
+ drout = -6.783373791e-01 ldrout = 3.008674840e-07 wdrout = 3.414318094e-12 pdrout = -8.510699994e-19
+ pscbe1 = 7.999049059e+08 lpscbe1 = 1.704715765e-02 wpscbe1 = 1.021465302e-06 ppscbe1 = -2.546157837e-13
+ pscbe2 = -6.326537659e-08 lpscbe2 = 1.797452289e-14 wpscbe2 = 5.923823942e-14 ppscbe2 = -1.476601975e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.042511144e+01 lbeta0 = -3.776776388e-07 wbeta0 = -6.630336816e-08 pbeta0 = 1.652710906e-14
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.848087777e-08 lagidl = -9.591657264e-15 wagidl = -2.987199179e-14 pagidl = 7.446042033e-21
+ bgidl = 1.854155595e+09 lbgidl = -1.531201946e+02 wbgidl = 3.791282654e-06 pbgidl = -9.450321198e-13
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.206339816e+00 lkt1 = 4.196324657e-07 wkt1 = 1.341456233e-06 pkt1 = -3.343780880e-13
+ kt2 = 1.609882469e+00 lkt2 = -4.144518324e-07 wkt2 = -1.211406378e-06 pkt2 = 3.019612108e-13
+ at = -6.479090521e+05 lat = 1.784230765e-01 wat = 6.121637171e-01 pat = -1.525909889e-7
+ ute = -1.762536546e+01 lute = 4.185353020e-06 wute = 1.154184163e-05 pute = -2.876977153e-12
+ ua1 = -1.428237563e-08 lua1 = 3.633638559e-15 wua1 = 1.048555150e-14 pua1 = -2.613680995e-21
+ ub1 = 1.284640297e-17 lub1 = -3.244364548e-24 wub1 = -9.556618169e-24 pub1 = 2.382130428e-30
+ uc1 = -5.435554732e-10 luc1 = 1.110897971e-16 wuc1 = 1.961246690e-16 puc1 = -4.888701562e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.143 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-9.691315548e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.765995610e-08 wvth0 = -5.784951806e-08 pvth0 = 2.155805425e-14
+ k1 = 3.789719604e+00 lk1 = -4.237772373e-07 wk1 = -2.030930521e-06 pk1 = 3.189421750e-13
+ k2 = -2.625016385e+00 lk2 = 3.911461170e-07 wk2 = 1.816263078e-06 pk2 = -2.963893501e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -8.220297122e+00 ldsub = 1.349322598e-06 wdsub = 6.466556141e-06 pdsub = -1.015523557e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {2.968393333e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.200469550e-07 wvoff = -2.491660809e-06 pvoff = 3.912695994e-13
+ nfactor = {2.542207029e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.449336086e-06 wnfactor = -1.652654432e-05 pnfactor = 2.595189714e-12
+ eta0 = -1.833050382e+01 leta0 = 2.934366908e-06 weta0 = 1.405920609e-05 peta0 = -2.207740225e-12
+ etab = -1.848093984e+00 letab = 2.880107474e-07 wetab = 1.380276236e-06 petab = -2.167618868e-13
+ u0 = 1.475278189e-01 lu0 = -2.283274774e-08 wu0 = -1.075382468e-07 pu0 = 1.711397984e-14
+ ua = 5.094477068e-08 lua = -8.300483604e-15 wua = -3.976946432e-14 pua = 6.245064782e-21
+ ub = -4.133425721e-17 lub = 6.775785315e-24 wub = 3.246430039e-23 pub = -5.097921860e-30
+ uc = 9.214243828e-10 luc = -1.457415584e-16 wuc = -6.984588321e-16 puc = 1.096876367e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.269448930e+05 lvsat = -8.600412034e-02 wvsat = -4.228705677e-01 pvsat = 6.581320991e-8
+ a0 = 1.869933686e+01 la0 = -2.778718950e-06 wa0 = -1.331346223e-05 pa0 = 2.090634713e-12
+ ags = 1.250000083e+00 lags = -1.372824698e-14 wags = -1.930405347e-14 pags = 3.209587263e-21
+ a1 = 0.0
+ a2 = -6.460558624e+00 la2 = 1.124022542e-06 wa2 = 5.386819554e-06 pa2 = -8.459589649e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.148466247e-01 lketa = -1.445944279e-07 wketa = -6.927839759e-07 pketa = 1.087890196e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.116745920e-01 lpclm = -1.417296317e-08 wpclm = -6.792328090e-08 ppclm = 1.066682322e-14
+ pdiblc1 = -1.269578008e+01 lpdiblc1 = 2.034809161e-06 wpdiblc1 = 9.751716875e-06 ppdiblc1 = -1.531432869e-12
+ pdiblc2 = 1.838890236e-01 lpdiblc2 = -2.847796511e-08 wpdiblc2 = -1.364791806e-07 ppdiblc2 = 2.143301445e-14
+ pdiblcb = 5.176138480e+01 lpdiblcb = -8.247913955e-06 wpdiblcb = -3.952769936e-05 ppdiblcb = 6.207523887e-12
+ drout = 1.000012181e+00 ldrout = -2.025304443e-12 wdrout = -8.722241716e-12 pdrout = 1.450203522e-18
+ pscbe1 = 8.000000041e+08 lpscbe1 = -6.799716949e-07 wpscbe1 = -2.609443665e-06 ppscbe1 = 4.338588715e-13
+ pscbe2 = 1.600607431e-07 lpscbe2 = -2.415202390e-14 wpscbe2 = -1.157473198e-13 ppscbe2 = 1.817723466e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.180557734e+00 lbeta0 = 2.703389157e-08 wbeta0 = 1.295561064e-07 pbeta0 = -2.034595729e-14
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -9.831766554e-08 lagidl = 1.634751593e-14 wagidl = 7.631645820e-14 pagidl = -1.268891348e-20
+ bgidl = 1.000000297e+09 lbgidl = -4.937791252e-05 wbgidl = -9.685241699e-06 pbgidl = 1.610313416e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.921126947e+00 lkt1 = -5.469153494e-07 wkt1 = -2.620393368e-06 pkt1 = 4.114846903e-13
+ kt2 = -3.218575971e+00 lkt2 = 4.939024023e-07 wkt2 = 2.367001600e-06 pkt2 = -3.717195439e-13
+ at = 1.619069260e+06 lat = -2.495852631e-01 wat = -1.196124390e+00 pat = 1.878422175e-7
+ ute = 2.969831120e+01 lute = -4.705724348e-06 wute = -2.255193939e-05 pute = 3.541610219e-12
+ ua1 = 2.776936883e-08 lua1 = -4.275063039e-15 wua1 = -2.048801836e-14 pua1 = 3.217486950e-21
+ ub1 = -2.510413376e-17 lub1 = 3.896329024e-24 wub1 = 1.867295362e-23 pub1 = -2.932445063e-30
+ uc1 = 4.835589388e-10 luc1 = -7.996198153e-17 wuc1 = -3.832136490e-16 puc1 = 6.018078184e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.144 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.145 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.120472155e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.870888723e-7
+ k1 = 4.170862753e-01 lk1 = 2.913759846e-7
+ k2 = 2.448249051e-02 lk2 = -5.836714509e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = 1.694065895e-27 pcit = 3.388131789e-32
+ voff = {-2.688785328e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.293878253e-7
+ nfactor = {2.183144685e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.000922662e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.113674562e-02 lu0 = -1.256245066e-8
+ ua = -9.216113352e-10 lua = 2.090566673e-15
+ ub = 1.520604476e-18 lub = -5.620003986e-24
+ uc = -1.046565291e-10 luc = -2.012847738e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.288282795e+04 lvsat = -2.545272048e-1
+ a0 = 1.626037978e+00 la0 = -3.240640463e-6
+ ags = 1.127453634e-01 lags = 1.089233216e-8
+ a1 = 0.0
+ a2 = 1.083322921e+00 la2 = -2.266375124e-6
+ b0 = -2.350169889e-07 lb0 = 2.106462362e-12
+ b1 = 4.206262362e-10 lb1 = 3.533945400e-15
+ keta = 3.418087999e-02 lketa = -2.163844674e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.896493835e-02 lpclm = 1.679237053e-06 wpclm = -2.775557562e-23 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.907724688e-03 lpdiblc2 = -1.261085430e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.864397580e-09 lpscbe2 = 2.392366917e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.666054167e-11 lalpha0 = 1.333161838e-15
+ alpha1 = -6.666054167e-11 lalpha1 = 1.333161838e-15
+ beta0 = 4.799834625e+01 lbeta0 = -3.599536962e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.809193870e-09 lagidl = -1.817806134e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443729441e-01 lkt1 = 1.224543810e-7
+ kt2 = -6.520326764e-02 lkt2 = 1.331404597e-07 wkt2 = 1.110223025e-22
+ at = 7.714160610e+04 lat = -1.230276006e-1
+ ute = 5.604140827e-01 lute = -1.286740876e-05 wute = -4.440892099e-22 pute = 7.105427358e-27
+ ua1 = 3.770448273e-09 lua1 = -3.360373048e-14
+ ub1 = -2.644626951e-18 lub1 = 2.831349847e-23 pub1 = 2.465190329e-44
+ uc1 = -9.425493132e-11 luc1 = 1.289271244e-15 wuc1 = -5.169878828e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.146 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.074934676e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.282250820e-8
+ k1 = 4.603687398e-01 lk1 = -5.485191820e-8
+ k2 = 1.663300362e-02 lk2 = 4.422980655e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.526831662e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.983679658e-08 wvoff = -4.440892099e-22
+ nfactor = {1.083406992e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.796170572e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.366897430e-03 lu0 = 9.594299004e-9
+ ua = -8.793373383e-10 lua = 1.752405770e-15
+ ub = 9.308044156e-19 lub = -9.020370027e-25
+ uc = -1.070081003e-10 luc = -1.317636748e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.342668478e+04 lvsat = -1.889970965e-2
+ a0 = 1.169514648e+00 la0 = 4.112106358e-7
+ ags = 4.518586659e-02 lags = 5.513186502e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.904470373e-08 lb0 = 7.415555649e-14
+ b1 = 2.692493660e-09 lb1 = -1.463932417e-14 pb1 = -6.617444900e-36
+ keta = 7.537928491e-03 lketa = -3.260437949e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.076066625e-01 lpclm = 4.388121945e-06 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 2.324642703e-04 lpdiblc2 = 7.899977302e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.461814170e-08 lpscbe2 = -2.210205481e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.999816250e-10 lalpha0 = -7.997795135e-16
+ alpha1 = 1.999816250e-10 lalpha1 = -7.997795135e-16
+ beta0 = -2.399503875e+01 lbeta0 = 2.159404686e-04 wbeta0 = -7.105427358e-21 pbeta0 = -2.842170943e-26
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.936827142e-10 lagidl = -1.255526991e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.138822703e-01 lkt1 = -1.214485986e-7
+ kt2 = -3.857419708e-02 lkt2 = -7.987253241e-8
+ at = 2.254069419e+04 lat = 3.137395630e-1
+ ute = -1.913180623e+00 lute = 6.919530795e-6
+ ua1 = -2.950544819e-09 lua1 = 2.015927433e-14 pua1 = -3.308722450e-36
+ ub1 = 2.918299229e-18 lub1 = -1.618582223e-23 wub1 = 3.081487911e-39
+ uc1 = 5.518884344e-10 luc1 = -3.879400767e-15 wuc1 = 2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.147 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.073354483e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.650289888e-8
+ k1 = 3.860761503e-01 lk1 = 2.422638348e-7
+ k2 = 3.864608706e-02 lk2 = -8.361317351e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.598897400e-01 ldsub = -1.199338541e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.344875018e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.706751263e-8
+ nfactor = {2.301599641e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.570464991e-8
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394744587e-01 letab = 2.778467713e-7
+ u0 = 1.198857651e-02 lu0 = -4.889755366e-9
+ ua = -1.319018025e-10 lua = -1.236787009e-15
+ ub = 5.490351914e-19 lub = 6.247592937e-25
+ uc = -1.334915649e-10 luc = 1.045967563e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.358762876e+04 lvsat = -9.952866729e-02 wvsat = 1.164153218e-16
+ a0 = 1.399225751e+00 la0 = -5.074649400e-7
+ ags = -4.159569572e-02 lags = 8.983811150e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.819412950e-08 lb0 = 7.755722824e-14
+ b1 = -2.575139163e-09 lb1 = 6.427335412e-15 pb1 = -6.617444900e-36
+ keta = 2.261809468e-02 lketa = -6.357001880e-08 pketa = 5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.069927487e-01 lpclm = 3.304700303e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.186804914e-04 lpdiblc2 = 4.526971437e-11
+ pdiblcb = -4.249265000e-01 lpdiblcb = 7.995590540e-07 wpdiblcb = -4.440892099e-22
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.717023012e-09 lpscbe2 = 1.498082628e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.996325000e-11 lalpha0 = 3.997795270e-16
+ alpha1 = -9.996325000e-11 lalpha1 = 3.997795270e-16
+ beta0 = 5.442312590e+01 lbeta0 = -9.767455261e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.805953197e-11 lagidl = 1.790882113e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.356331678e-01 lkt1 = -3.446099523e-8
+ kt2 = -6.315530546e-02 lkt2 = 1.843383399e-8
+ at = 1.619156016e+05 lat = -2.436576261e-1
+ ute = -9.264321097e-02 lute = -3.612807586e-7
+ ua1 = 2.877410594e-09 lua1 = -3.148263775e-15
+ ub1 = -1.895518164e-18 lub1 = 3.065909193e-24
+ uc1 = -8.716392777e-10 luc1 = 1.813663789e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.148 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.086028606e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.184182979e-8
+ k1 = 5.064839054e-01 lk1 = 1.536824197e-9
+ k2 = -2.175514322e-03 lk2 = -1.999974616e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000200e-01 ldsub = -1.997795618e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.136546851e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.458280866e-8
+ nfactor = {2.242862352e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.172675677e-8
+ eta0 = -4.886402175e-01 leta0 = 9.779209169e-07 weta0 = 2.602085214e-23 peta0 = -7.979727989e-29
+ etab = 2.464242746e-04 letab = -1.492299927e-9
+ u0 = 1.041902600e-02 lu0 = -1.751807974e-9
+ ua = -6.756220924e-10 lua = -1.497460633e-16
+ ub = 8.575638770e-19 lub = 7.928691116e-27
+ uc = -1.187352451e-10 luc = 7.509496275e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.581072052e+04 lvsat = 3.597533316e-2
+ a0 = 1.033650996e+00 la0 = 2.234158726e-7
+ ags = 2.513648550e-01 lags = 3.126753396e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 8.083645775e-08 lb0 = -4.768138616e-14 wb0 = 1.058791184e-28
+ b1 = 4.795263422e-09 lb1 = -8.308052512e-15 wb1 = -1.654361225e-30 pb1 = 3.308722450e-36
+ keta = -1.731434613e-02 lketa = 1.626551248e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.164189562e-01 lpclm = -2.881549565e-7
+ pdiblc1 = 3.956566993e-01 lpdiblc1 = -1.130924086e-8
+ pdiblc2 = 4.526390171e-04 lpdiblc2 = -2.262237742e-11
+ pdiblcb = 1.748530000e-01 lpdiblcb = -3.995591080e-7
+ drout = 3.837641586e-01 ldrout = 3.523421494e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.762341479e-09 lpscbe2 = -5.917859960e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.665153203e+00 lbeta0 = 1.804820678e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.216142405e-10 lagidl = 8.118944782e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.266945131e-01 lkt1 = -5.233173475e-8
+ kt2 = -5.930686777e-02 lkt2 = 1.073978722e-8
+ at = 2.833087101e+04 lat = 2.341365030e-2
+ ute = 5.008903148e-01 lute = -1.547911563e-06 pute = 8.881784197e-28
+ ua1 = 3.034530159e-09 lua1 = -3.462387422e-15
+ ub1 = -1.577991139e-18 lub1 = 2.431088525e-24 wub1 = -7.703719778e-40 pub1 = -7.703719778e-46
+ uc1 = 4.156291695e-12 luc1 = 6.271635987e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.149 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.096247150e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.205286336e-08 wvth0 = 1.984942204e-08 pvth0 = -1.983483272e-14
+ k1 = -3.231479595e-01 lk1 = 8.305589096e-07 wk1 = 6.024375721e-07 pk1 = -6.019947805e-13
+ k2 = 3.416021413e-01 lk2 = -3.455249536e-07 wk2 = -2.524438723e-07 pk2 = 2.522583261e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.743818839e+00 ldsub = -7.478318232e-06 wdsub = -5.478904364e-06 pdsub = 5.474877369e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-5.861139759e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.576027246e-07 wvoff = 2.451297270e-07 pvoff = -2.449495566e-13
+ nfactor = {1.680825599e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.451296131e-05 wnfactor = -1.039972865e-05 pnfactor = 1.039208485e-11
+ eta0 = -4.401373598e+00 leta0 = 4.887778438e-06 weta0 = 3.579757738e-06 peta0 = -3.577126616e-12
+ etab = -5.674885495e-03 letab = 4.424657680e-09 wetab = 2.786050950e-09 petab = -2.784003203e-15
+ u0 = 7.431856396e-02 lu0 = -6.560437977e-08 wu0 = -4.621124007e-08 pu0 = 4.617727481e-14
+ ua = 6.864089159e-09 lua = -7.683915627e-15 wua = -5.312963977e-15 pua = 5.309058948e-21
+ ub = 3.226633454e-18 lub = -2.359399620e-24 wub = -1.983747723e-24 pub = 1.982289668e-30
+ uc = -2.462765338e-10 luc = 2.025425085e-16 wuc = 1.382144101e-16 puc = -1.381128225e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.044894211e+05 lvsat = 6.558195542e-01 wvsat = 4.296681730e-01 pvsat = -4.293523669e-7
+ a0 = 5.835613232e+00 la0 = -4.575016922e-06 wa0 = -2.955534113e-06 pa0 = 2.953361796e-12
+ ags = -1.204516165e-01 lags = 6.842185259e-07 wags = -4.757492178e-16 pags = 4.754010519e-22
+ a1 = 0.0
+ a2 = -4.444669312e+00 la2 = 5.240814480e-06 wa2 = 3.699404703e-06 pa2 = -3.696685641e-12
+ b0 = 6.619131254e-08 lb0 = -3.304700513e-14 wb0 = 7.063939260e-22 pb0 = -7.058747478e-28
+ b1 = -7.032627217e-09 lb1 = 3.511144628e-15 wb1 = 2.936822047e-25 pb1 = -2.934638290e-31
+ keta = -2.342131666e-02 lketa = 2.236799439e-08 wketa = 4.318775248e-08 pketa = -4.315600948e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.335355382e+00 lpclm = -4.703843464e-06 wpclm = -3.006429817e-06 ppclm = 3.004220091e-12
+ pdiblc1 = 1.354778486e+00 lpdiblc1 = -9.697260727e-07 wpdiblc1 = -4.373903697e-07 ppdiblc1 = 4.370688878e-13
+ pdiblc2 = 8.570039306e-03 lpdiblc2 = -8.134056378e-09 wpdiblc2 = -5.672394280e-09 ppdiblc2 = 5.668225070e-15
+ pdiblcb = -2.516041031e+00 lpdiblcb = 2.289357116e-06 wpdiblcb = 1.526548132e-06 ppdiblcb = -1.525426119e-12
+ drout = -4.481149613e+00 ldrout = 5.213680210e-06 wdrout = 3.625787154e-06 pdrout = -3.623122200e-12
+ pscbe1 = -5.917514882e+09 lpscbe1 = 6.712577509e+03 wpscbe1 = 4.916221465e+03 ppscbe1 = -4.912608042e-3
+ pscbe2 = 7.079213409e-07 lpscbe2 = -6.982376385e-13 wpscbe2 = -5.114974182e-13 ppscbe2 = 5.111214676e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.052914264e+00 lbeta0 = 5.414404622e-06 wbeta0 = 2.299086262e-06 pbeta0 = -2.297396434e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.259494204e-08 lagidl = -1.135248592e-14 wagidl = -7.356483322e-15 pagidl = 7.351076307e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.299727628e-01 lkt1 = -6.085898602e-07 wkt1 = -4.026052475e-07 pkt1 = 4.023093326e-13
+ kt2 = -3.372967282e-01 lkt2 = 2.885253251e-07 wkt2 = 1.996978499e-07 pkt2 = -1.995510720e-13
+ at = 5.243093137e+05 lat = -4.722002482e-01 wat = -3.336519476e-01 pat = 3.334067135e-7
+ ute = -2.303095054e+00 lute = 1.254012877e-06 wute = 2.975519563e-07 pute = -2.973332556e-13
+ ua1 = -1.256854174e-08 lua1 = 1.212921622e-14 wua1 = 6.693247224e-15 pua1 = -6.688327687e-21
+ ub1 = 2.010357870e-17 lub1 = -1.923454537e-23 wub1 = -1.168038137e-23 pub1 = 1.167179628e-29
+ uc1 = 1.628002898e-09 luc1 = -1.559936719e-15 wuc1 = -9.508363578e-16 puc1 = 9.501374930e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.150 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.483861333e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.176896731e-08 wvth0 = -3.969884408e-08 pvth0 = 9.895532370e-15
+ k1 = 2.100724792e+00 lk1 = -3.795959195e-07 wk1 = -1.204875144e-06 pk1 = 3.003332028e-13
+ k2 = -6.835814912e-01 lk2 = 1.663133526e-07 wk2 = 5.048877447e-07 pk2 = -1.258508437e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.523068623e+01 ldsub = 3.992048042e-06 wdsub = 1.095780873e-05 pdsub = -2.731398192e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {5.006193357e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.849651822e-07 wvoff = -4.902594540e-07 pvoff = 1.222045228e-13
+ nfactor = {-2.714331223e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.430518394e-06 wnfactor = 2.079945730e-05 pnfactor = -5.184576724e-12
+ eta0 = 1.027274719e+01 leta0 = -2.438496479e-06 weta0 = -7.159515476e-06 peta0 = 1.784616625e-12
+ etab = 6.437137313e-03 letab = -1.622451387e-09 wetab = -5.572101901e-09 petab = 1.388929980e-15
+ u0 = -1.208286600e-01 lu0 = 3.182579899e-08 wu0 = 9.242248013e-08 pu0 = -2.303768951e-14
+ ua = -1.572728623e-08 lua = 3.595167408e-15 wua = 1.062592795e-14 pua = -2.648671931e-21
+ ub = -4.577934267e-18 lub = 1.537147884e-24 wub = 3.967495445e-24 pub = -9.889577521e-31
+ uc = 3.193279093e-10 luc = -7.984399375e-17 wuc = -2.764288202e-16 puc = 6.890402988e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.317882333e+06 lvsat = -3.039533794e-01 wvsat = -8.593363459e-01 pvsat = 2.142024743e-7
+ a0 = -7.259650523e+00 la0 = 1.962989937e-06 wa0 = 5.911068226e-06 pa0 = -1.473422421e-12
+ ags = 9.950076816e-01 lags = 1.273087395e-07 wags = 9.514984356e-16 pags = -2.371747243e-22
+ a1 = 0.0
+ a2 = 1.129330499e+01 la2 = -2.616605258e-06 wa2 = -7.398809407e-06 pa2 = 1.844264227e-12
+ b0 = 2.120309864e-15 lb0 = -5.285190384e-22 wb0 = -1.412787906e-21 pb0 = 3.521585775e-28
+ b1 = 8.815098761e-19 lb1 = -2.197295593e-25 wb1 = -5.873606086e-25 pb1 = 1.464084421e-31
+ keta = 7.428292398e-02 lketa = -2.641231331e-08 wketa = -8.637550496e-08 pketa = 2.153039024e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -8.795676865e+00 lpclm = 2.351286351e-06 wpclm = 6.012859634e-06 ppclm = -1.498795457e-12
+ pdiblc1 = -1.576770556e+00 lpdiblc1 = 4.938937598e-07 wpdiblc1 = 8.747807394e-07 ppdiblc1 = -2.180522210e-13
+ pdiblc2 = -2.397263968e-02 lpdiblc2 = 8.113364246e-09 wpdiblc2 = 1.134478856e-08 ppdiblc2 = -2.827858720e-15
+ pdiblcb = 4.419916636e+00 lpdiblcb = -1.173523789e-06 wpdiblcb = -3.053096263e-06 ppdiblcb = 7.610300401e-13
+ drout = 1.137846932e+01 ldrout = -2.704472439e-06 wdrout = -7.251574308e-06 pdrout = 1.807563670e-12
+ pscbe1 = 1.423505639e+10 lpscbe1 = -3.348895988e+03 wpscbe1 = -9.832442931e+03 ppscbe1 = 2.450883887e-3
+ pscbe2 = -1.388007876e-06 lpscbe2 = 3.481864621e-13 wpscbe2 = 1.022994836e-12 ppscbe2 = -2.549968079e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.487660039e+01 lbeta0 = -1.487278032e-06 wbeta0 = -4.598172524e-06 pbeta0 = 1.146163474e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.025820368e-08 lagidl = 5.049939874e-15 wagidl = 1.471296664e-14 pagidl = -3.667427630e-21
+ bgidl = 7.608364006e+08 lbgidl = 1.194060145e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.653472721e+00 lkt1 = 2.818220495e-07 wkt1 = 8.052104950e-07 pkt1 = -2.007107940e-13
+ kt2 = 5.331574119e-01 lkt2 = -1.460619611e-07 wkt2 = -3.993956998e-07 pkt2 = 9.955536910e-14
+ at = -9.094119413e+05 lat = 2.436065941e-01 wat = 6.673038953e-01 pat = -1.663355055e-7
+ ute = 1.248767304e+00 lute = -5.193076834e-07 wute = -5.951039125e-07 pute = 1.483385768e-13
+ ua1 = 2.312256412e-08 lua1 = -5.690103746e-15 wua1 = -1.338649445e-14 pua1 = 3.336784539e-21
+ ub1 = -3.662130493e-17 lub1 = 9.086203661e-24 wub1 = 2.336076273e-23 pub1 = -5.823020522e-30
+ uc1 = -2.890929178e-09 luc1 = 6.962079037e-16 wuc1 = 1.901672716e-15 puc1 = -4.740204494e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.151 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.981652160e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.428728428e-8
+ k1 = -6.868110801e-01 lk1 = 3.152392096e-7
+ k2 = 4.810608589e-01 lk2 = -1.239912228e-07 wk2 = 2.220446049e-22 pk2 = 9.714451465e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.682474392e+00 ldsub = -2.238109408e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {8.041300560e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.022245136e-8
+ nfactor = {1.047285534e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.035890417e-7
+ eta0 = 4.900000008e-01 leta0 = -5.696065841e-17
+ etab = 1.925516612e-03 letab = -4.978622536e-10 wetab = 8.673617380e-25 petab = 5.421010862e-32
+ u0 = 1.623006395e-02 lu0 = -2.338143833e-9
+ ua = 1.228104028e-09 lua = -6.312179456e-16
+ ub = 2.170685950e-19 lub = 3.419214952e-25
+ uc = 3.061872191e-11 luc = -7.878898151e-18 wuc = -6.462348536e-33 puc = -8.077935669e-40
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.760102185e+05 lvsat = -1.932462687e-2
+ a0 = -5.465138832e-02 la0 = 1.670358279e-7
+ ags = 2.160686824e+00 lags = -1.632542721e-7
+ a1 = 0.0
+ a2 = 9.172257814e-01 la2 = -3.021187522e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.064756593e-02 lketa = 1.220643526e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.792752505e-01 lpclm = -1.048758818e-8
+ pdiblc1 = 5.315421921e-01 lpdiblc1 = -3.163481747e-8
+ pdiblc2 = 2.737215973e-02 lpdiblc2 = -4.685097180e-9
+ pdiblcb = 1.891439592e+00 lpdiblcb = -5.432629582e-7
+ drout = -6.783326782e-01 ldrout = 3.008663122e-7
+ pscbe1 = 7.999049073e+08 lpscbe1 = 1.704680709e-2
+ pscbe2 = 1.829494379e-08 lpscbe2 = -2.355610367e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.033382372e+01 lbeta0 = -3.549228047e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.647441449e-09 lagidl = 6.601932258e-16 wagidl = -1.479877815e-30 pagidl = 2.488004186e-37
+ bgidl = 1.854155600e+09 lbgidl = -1.531201959e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.593976841e-01 lkt1 = -4.074556472e-8
+ kt2 = -5.800457968e-02 lkt2 = 1.294032692e-9
+ at = 1.949294486e+05 lat = -3.166706240e-02 wat = -2.328306437e-16
+ ute = -1.734341181e+00 lute = 2.242768531e-7
+ ua1 = 1.543285759e-10 lua1 = 3.507348664e-17
+ ub1 = -3.113283727e-19 lub1 = 3.539735529e-26
+ uc1 = -2.735273461e-10 luc1 = 4.378123603e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.152 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-5.973392663e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.658040985e-08 wvth0 = -3.278867187e-07 pvth0 = 6.435268685e-14
+ k1 = 1.250497272e-01 lk1 = 1.857940101e-07 wk1 = 6.307631871e-07 pk1 = -1.237967369e-13
+ k2 = 8.334985177e-01 lk2 = -2.049206951e-07 wk2 = -6.956977978e-07 pk2 = 1.365411283e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.448137155e+00 ldsub = -5.915731091e-07 wdsub = -2.008367695e-06 pdsub = 3.941722857e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.518026053e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.258875611e-07 wvoff = 7.668794275e-07 pvoff = -1.505115908e-13
+ nfactor = {-4.335228634e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.498261209e-06 wnfactor = 5.086538978e-06 pnfactor = -9.983095726e-13
+ eta0 = 6.984138676e+00 leta0 = -1.274572127e-06 weta0 = -4.327122528e-06 peta0 = 8.492627029e-13
+ etab = 6.425158375e-01 letab = -1.262705347e-07 wetab = -4.286835647e-07 petab = 8.413557983e-14
+ u0 = -4.184376791e-02 lu0 = 8.837986683e-09 wu0 = 3.000460916e-08 pu0 = -5.888854617e-15
+ ua = -2.066308686e-08 lua = 3.605397180e-15 wua = 1.224018191e-14 pua = -2.402319302e-21
+ ub = 1.712008569e-17 lub = -2.943124167e-24 wub = -9.991790301e-24 pub = 1.961038723e-30
+ uc = -3.388951992e-10 luc = 6.389658248e-17 wuc = 2.169264041e-16 puc = -4.257506070e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.160462853e+05 lvsat = 5.578975612e-02 wvsat = 1.894040409e-01 pvsat = -3.717338409e-8
+ a0 = -5.272543711e+00 la0 = 1.206965752e-06 wa0 = 4.097602297e-06 pa0 = -8.042159147e-13
+ ags = 1.250000055e+00 lags = -9.178648952e-15 wags = 4.832401146e-16 pags = -9.484146801e-23
+ a1 = 0.0
+ a2 = 3.259576106e+00 la2 = -4.927983043e-07 wa2 = -1.673030942e-06 pa2 = 3.283574178e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.325616248e-01 lketa = 6.280590470e-08 wketa = 2.132236046e-07 pketa = -4.184833077e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.891113482e-01 lpclm = 6.213874579e-09 wpclm = 2.109587385e-08 ppclm = -4.140381681e-15
+ pdiblc1 = 4.900501202e+00 lpdiblc1 = -8.921085402e-07 wpdiblc1 = -3.028673379e-06 ppdiblc1 = 5.944225806e-13
+ pdiblc2 = -6.237804465e-02 lpdiblc2 = 1.248543108e-08 wpdiblc2 = 4.238754622e-08 ppdiblc2 = -8.319191760e-15
+ pdiblcb = -1.956355689e+01 lpdiblcb = 3.616083391e-06 wpdiblcb = 1.227646169e-05 ppdiblcb = -2.409439753e-12
+ drout = 1.000000198e+00 ldrout = -3.384324287e-14 wdrout = -1.926657234e-14 pdrout = 3.781353897e-21
+ pscbe1 = 8.000000016e+08 lpscbe1 = -3.117389679e-07 wpscbe1 = -8.478698730e-07 ppscbe1 = 1.664066315e-13
+ pscbe2 = -4.879710325e-08 lpscbe2 = 1.058882377e-14 wpscbe2 = 3.594864032e-14 ppscbe2 = -7.055459893e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.414325248e+00 lbeta0 = -1.185036134e-08 wbeta0 = -4.023204450e-08 pbeta0 = 7.896142215e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 7.028836208e-08 lagidl = -1.359194502e-14 wagidl = -4.614412293e-14 pagidl = 9.056476287e-21
+ bgidl = 1.000000267e+09 lbgidl = -4.383736801e-05 wbgidl = 1.229892731e-05 pbgidl = -2.413848877e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.797083967e+00 lkt1 = 2.375579635e-07 wkt1 = 8.064998375e-07 pkt1 = -1.582876906e-13
+ kt2 = 1.052511930e+00 lkt2 = -2.165387749e-07 wkt2 = -7.351407963e-07 pkt2 = 1.442824084e-13
+ at = -5.392527451e+05 lat = 1.094241653e-01 wat = 3.714907827e-01 pat = -7.291063846e-8
+ ute = -1.099506875e+01 lute = 2.063102099e-06 wute = 7.004150796e-06 pute = -1.374669656e-12
+ ua1 = -9.199820866e-09 lua1 = 1.874291704e-15 wua1 = 6.363147744e-15 pua1 = -1.248863192e-21
+ ub1 = 8.589890721e-18 lub1 = -1.708243620e-24 wub1 = -5.799420697e-24 pub1 = 1.138223303e-30
+ uc1 = -2.079230570e-10 luc1 = 3.505725813e-17 wuc1 = 1.190180224e-16 puc1 = -2.335907216e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.153 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.154 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.120472155e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.870888723e-7
+ k1 = 4.170862753e-01 lk1 = 2.913759846e-7
+ k2 = 2.448249051e-02 lk2 = -5.836714509e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = -2.371692252e-26 pcit = 3.523657061e-31
+ voff = {-2.688785328e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.293878253e-7
+ nfactor = {2.183144685e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.000922662e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.113674562e-02 lu0 = -1.256245066e-8
+ ua = -9.216113352e-10 lua = 2.090566673e-15
+ ub = 1.520604476e-18 lub = -5.620003986e-24
+ uc = -1.046565291e-10 luc = -2.012847738e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.288282795e+04 lvsat = -2.545272048e-1
+ a0 = 1.626037978e+00 la0 = -3.240640463e-6
+ ags = 1.127453634e-01 lags = 1.089233216e-8
+ a1 = 0.0
+ a2 = 1.083322921e+00 la2 = -2.266375124e-6
+ b0 = -2.350169889e-07 lb0 = 2.106462362e-12
+ b1 = 4.206262362e-10 lb1 = 3.533945400e-15
+ keta = 3.418087999e-02 lketa = -2.163844674e-07 pketa = -1.776356839e-27
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.896493835e-02 lpclm = 1.679237053e-06 wpclm = 2.220446049e-22 ppclm = -7.105427358e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.907724688e-03 lpdiblc2 = -1.261085430e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.864397580e-09 lpscbe2 = 2.392366917e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.666054167e-11 lalpha0 = 1.333161838e-15
+ alpha1 = -6.666054167e-11 lalpha1 = 1.333161838e-15
+ beta0 = 4.799834625e+01 lbeta0 = -3.599536962e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.809193870e-09 lagidl = -1.817806134e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443729441e-01 lkt1 = 1.224543810e-7
+ kt2 = -6.520326764e-02 lkt2 = 1.331404597e-7
+ at = 7.714160610e+04 lat = -1.230276006e-1
+ ute = 5.604140827e-01 lute = -1.286740876e-05 wute = 8.881784197e-22 pute = -2.842170943e-26
+ ua1 = 3.770448273e-09 lua1 = -3.360373048e-14 wua1 = -2.646977960e-29
+ ub1 = -2.644626951e-18 lub1 = 2.831349847e-23
+ uc1 = -9.425493132e-11 luc1 = 1.289271244e-15 wuc1 = -4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.155 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.074934676e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.282250820e-8
+ k1 = 4.603687398e-01 lk1 = -5.485191820e-8
+ k2 = 1.663300362e-02 lk2 = 4.422980655e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.526831662e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.983679658e-8
+ nfactor = {1.083406992e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.796170572e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.366897430e-03 lu0 = 9.594299004e-9
+ ua = -8.793373383e-10 lua = 1.752405770e-15 wua = 6.617444900e-30
+ ub = 9.308044156e-19 lub = -9.020370027e-25
+ uc = -1.070081003e-10 luc = -1.317636749e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.342668478e+04 lvsat = -1.889970965e-2
+ a0 = 1.169514648e+00 la0 = 4.112106358e-7
+ ags = 4.518586659e-02 lags = 5.513186502e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.904470373e-08 lb0 = 7.415555649e-14
+ b1 = 2.692493660e-09 lb1 = -1.463932417e-14
+ keta = 7.537928491e-03 lketa = -3.260437949e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.076066625e-01 lpclm = 4.388121945e-06 wpclm = 1.776356839e-21 ppclm = 7.105427358e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 2.324642703e-04 lpdiblc2 = 7.899977302e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.461814170e-08 lpscbe2 = -2.210205481e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.999816250e-10 lalpha0 = -7.997795135e-16
+ alpha1 = 1.999816250e-10 lalpha1 = -7.997795135e-16
+ beta0 = -2.399503875e+01 lbeta0 = 2.159404686e-04 pbeta0 = -2.273736754e-25
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.936827142e-10 lagidl = -1.255526991e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.138822703e-01 lkt1 = -1.214485986e-7
+ kt2 = -3.857419708e-02 lkt2 = -7.987253241e-8
+ at = 2.254069419e+04 lat = 3.137395630e-1
+ ute = -1.913180623e+00 lute = 6.919530795e-6
+ ua1 = -2.950544819e-09 lua1 = 2.015927433e-14 wua1 = -1.323488980e-29
+ ub1 = 2.918299229e-18 lub1 = -1.618582223e-23
+ uc1 = 5.518884344e-10 luc1 = -3.879400767e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.156 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.073354483e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.650289887e-8
+ k1 = 3.860761503e-01 lk1 = 2.422638348e-7
+ k2 = 3.864608706e-02 lk2 = -8.361317351e-08 wk2 = -2.220446049e-22
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.598897400e-01 ldsub = -1.199338541e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.344875018e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.706751263e-8
+ nfactor = {2.301599641e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.570464991e-8
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394744587e-01 letab = 2.778467713e-7
+ u0 = 1.198857651e-02 lu0 = -4.889755366e-9
+ ua = -1.319018025e-10 lua = -1.236787009e-15
+ ub = 5.490351914e-19 lub = 6.247592937e-25
+ uc = -1.334915649e-10 luc = 1.045967563e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.358762876e+04 lvsat = -9.952866729e-2
+ a0 = 1.399225751e+00 la0 = -5.074649400e-7
+ ags = -4.159569572e-02 lags = 8.983811150e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.819412950e-08 lb0 = 7.755722824e-14
+ b1 = -2.575139163e-09 lb1 = 6.427335412e-15 pb1 = -2.646977960e-35
+ keta = 2.261809468e-02 lketa = -6.357001880e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.069927487e-01 lpclm = 3.304700303e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.186804914e-04 lpdiblc2 = 4.526971437e-11
+ pdiblcb = -4.249265000e-01 lpdiblcb = 7.995590540e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.717023012e-09 lpscbe2 = 1.498082628e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.996325000e-11 lalpha0 = 3.997795270e-16
+ alpha1 = -9.996325000e-11 lalpha1 = 3.997795270e-16
+ beta0 = 5.442312590e+01 lbeta0 = -9.767455261e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.805953197e-11 lagidl = 1.790882113e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.356331678e-01 lkt1 = -3.446099523e-8
+ kt2 = -6.315530546e-02 lkt2 = 1.843383399e-8
+ at = 1.619156016e+05 lat = -2.436576261e-1
+ ute = -9.264321097e-02 lute = -3.612807586e-7
+ ua1 = 2.877410594e-09 lua1 = -3.148263775e-15
+ ub1 = -1.895518164e-18 lub1 = 3.065909193e-24
+ uc1 = -8.716392777e-10 luc1 = 1.813663789e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.157 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.086028606e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.184182979e-8
+ k1 = 5.064839054e-01 lk1 = 1.536824197e-9
+ k2 = -2.175514322e-03 lk2 = -1.999974616e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000200e-01 ldsub = -1.997796062e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.136546851e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.458280866e-8
+ nfactor = {2.242862352e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.172675677e-8
+ eta0 = -4.886402175e-01 leta0 = 9.779209169e-07 weta0 = -2.706168623e-22 peta0 = 2.768618668e-27
+ etab = 2.464242746e-04 letab = -1.492299927e-09 petab = 6.938893904e-30
+ u0 = 1.041902600e-02 lu0 = -1.751807974e-9
+ ua = -6.756220924e-10 lua = -1.497460633e-16
+ ub = 8.575638770e-19 lub = 7.928691116e-27
+ uc = -1.187352451e-10 luc = 7.509496275e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.581072052e+04 lvsat = 3.597533316e-2
+ a0 = 1.033650996e+00 la0 = 2.234158726e-7
+ ags = 2.513648550e-01 lags = 3.126753396e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 8.083645776e-08 lb0 = -4.768138616e-14
+ b1 = 4.795263422e-09 lb1 = -8.308052512e-15 wb1 = -1.323488980e-29 pb1 = 6.617444900e-36
+ keta = -1.731434613e-02 lketa = 1.626551248e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.164189562e-01 lpclm = -2.881549565e-7
+ pdiblc1 = 3.956566993e-01 lpdiblc1 = -1.130924086e-8
+ pdiblc2 = 4.526390171e-04 lpdiblc2 = -2.262237742e-11
+ pdiblcb = 1.748530000e-01 lpdiblcb = -3.995591080e-07 wpdiblcb = -4.440892099e-22
+ drout = 3.837641586e-01 ldrout = 3.523421494e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.762341479e-09 lpscbe2 = -5.917859960e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.665153203e+00 lbeta0 = 1.804820678e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.216142405e-10 lagidl = 8.118944782e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.266945131e-01 lkt1 = -5.233173475e-8
+ kt2 = -5.930686777e-02 lkt2 = 1.073978722e-8
+ at = 2.833087101e+04 lat = 2.341365030e-2
+ ute = 5.008903148e-01 lute = -1.547911563e-06 pute = 3.552713679e-27
+ ua1 = 3.034530159e-09 lua1 = -3.462387422e-15 wua1 = -1.323488980e-29
+ ub1 = -1.577991139e-18 lub1 = 2.431088525e-24
+ uc1 = 4.156291695e-12 luc1 = 6.271635987e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.158 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.066457169e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.228477766e-8
+ k1 = 5.809893998e-01 lk1 = -7.291390867e-8
+ k2 = -3.726522465e-02 lk2 = 3.306394477e-08 wk2 = 5.551115123e-23 pk2 = -5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.789122000e-01 ldsub = 7.383690995e-07 pdsub = -1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.182236678e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.001718417e-8
+ nfactor = {1.200359609e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.083463260e-6
+ eta0 = 9.711211764e-01 leta0 = -4.807675523e-7
+ etab = -1.493584618e-03 letab = 2.464300584e-10
+ u0 = 4.964807659e-03 lu0 = 3.698401517e-9
+ ua = -1.109598808e-09 lua = 2.839116794e-16
+ ub = 2.494279967e-19 lub = 6.156175915e-25
+ uc = -3.884456477e-11 luc = -4.736997978e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.035589602e+04 lvsat = 1.144819836e-2
+ a0 = 1.399952291e+00 la0 = -1.426161911e-7
+ ags = -1.204516172e-01 lags = 6.842185266e-7
+ a1 = 0.0
+ a2 = 1.107391439e+00 la2 = -3.071655067e-7
+ b0 = 6.619131360e-08 lb0 = -3.304700618e-14
+ b1 = -7.032627217e-09 lb1 = 3.511144627e-15
+ keta = 4.139479423e-02 lketa = -4.240047666e-08 wketa = -4.163336342e-23
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.233102479e-01 lpclm = -1.951146831e-7
+ pdiblc1 = 6.983437078e-01 lpdiblc1 = -3.137737744e-7
+ pdiblc2 = 5.691890659e-05 lpdiblc2 = 3.728068788e-10
+ pdiblcb = -0.225
+ drout = 9.604260361e-01 ldrout = -2.238958816e-7
+ pscbe1 = 1.460742549e+09 lpscbe1 = -6.602569028e+2
+ pscbe2 = -5.973317864e-08 lpscbe2 = 6.885265491e-14 wpscbe2 = -2.117582368e-28 ppscbe2 = -2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.503379304e+00 lbeta0 = 1.966475673e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.554343458e-09 lagidl = -3.200021832e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.742565584e-01 lkt1 = -4.804647554e-9
+ kt2 = -3.759050968e-02 lkt2 = -1.096060934e-8
+ at = 2.356499624e+04 lat = 2.817602215e-2
+ ute = -1.856529547e+00 lute = 8.077755953e-07 pute = 7.105427358e-27
+ ua1 = -2.523326854e-09 lua1 = 2.091384566e-15
+ ub1 = 2.573680751e-18 lub1 = -1.717531887e-24 wub1 = 1.232595164e-38 pub1 = -6.162975822e-45
+ uc1 = 2.009891904e-10 luc1 = -1.339718666e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.159 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.007966096e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.917767921e-9
+ k1 = 2.924500733e-01 lk1 = 7.114367819e-8
+ k2 = 7.415324063e-02 lk2 = -2.256339530e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.214775846e+00 ldsub = -1.072300629e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.351612806e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.560826904e-9
+ nfactor = {4.072480519e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.504861863e-7
+ eta0 = -4.722423533e-01 leta0 = 2.398533403e-07 weta0 = -1.776356839e-21 peta0 = -3.053113318e-28
+ etab = -1.925464442e-03 letab = 4.620525390e-10
+ u0 = 1.787885262e-02 lu0 = -2.749129141e-9
+ ua = 2.200897025e-10 lua = -3.799552548e-16
+ ub = 1.376476647e-18 lub = 5.292164706e-26
+ uc = -9.553602869e-11 luc = 2.356706576e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.819169822e+04 lvsat = 1.752135658e-2
+ a0 = 1.611671360e+00 la0 = -2.483201119e-7
+ ags = 9.950076830e-01 lags = 1.273087391e-7
+ a1 = 0.0
+ a2 = 1.891834845e-01 la2 = 1.512635879e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.534929780e-02 lketa = 5.900462451e-09 wketa = -4.440892099e-22
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.284134026e-01 lpclm = 1.018964903e-7
+ pdiblc1 = -2.639010008e-01 lpdiblc1 = 1.666413300e-07 wpdiblc1 = -8.881784197e-22
+ pdiblc2 = -6.946398880e-03 lpdiblc2 = 3.869318333e-09 wpdiblc2 = 1.387778781e-23 ppdiblc2 = 1.387778781e-29
+ pdiblcb = -1.621654265e-01 lpdiblcb = -3.137110336e-8
+ drout = 4.953180247e-01 ldrout = 8.316269749e-9
+ pscbe1 = -5.214584712e+08 lpscbe1 = 3.293866893e+02 wpscbe1 = 1.907348633e-12 ppscbe1 = 4.768371582e-19
+ pscbe2 = 1.473011627e-07 lpscbe2 = -3.451234553e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.975670309e+00 lbeta0 = 2.328823045e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.822993481e-09 lagidl = -4.541297369e-16
+ bgidl = 7.608364006e+08 lbgidl = 1.194060145e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.450140790e-01 lkt1 = -1.940439406e-8
+ kt2 = -6.625502520e-02 lkt2 = 3.350579994e-9
+ at = 9.207669362e+04 lat = -6.029470441e-3
+ ute = 3.556362895e-01 lute = -2.966813811e-07 pute = -8.881784197e-28
+ ua1 = 3.032134340e-09 lua1 = -6.822627670e-16
+ ub1 = -1.561509020e-18 lub1 = 3.470236344e-25
+ uc1 = -3.690176234e-11 luc1 = -1.520124011e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.160 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.981652160e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.428728428e-8
+ k1 = -6.868110801e-01 lk1 = 3.152392096e-7
+ k2 = 4.810608589e-01 lk2 = -1.239912228e-07 wk2 = 8.881784197e-22 pk2 = -2.220446049e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.682474392e+00 ldsub = -2.238109408e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {8.041300560e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.022245136e-8
+ nfactor = {1.047285534e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.035890417e-7
+ eta0 = 4.900000008e-01 leta0 = -5.696065841e-17
+ etab = 1.925516612e-03 letab = -4.978622536e-10 wetab = 6.938893904e-24 petab = 1.734723476e-30
+ u0 = 1.623006395e-02 lu0 = -2.338143833e-9
+ ua = 1.228104028e-09 lua = -6.312179456e-16
+ ub = 2.170685950e-19 lub = 3.419214952e-25
+ uc = 3.061872191e-11 luc = -7.878898151e-18 wuc = -5.169878828e-32 puc = 2.584939414e-38
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.760102185e+05 lvsat = -1.932462687e-2
+ a0 = -5.465138832e-02 la0 = 1.670358279e-7
+ ags = 2.160686824e+00 lags = -1.632542721e-7
+ a1 = 0.0
+ a2 = 9.172257814e-01 la2 = -3.021187522e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.064756593e-02 lketa = 1.220643526e-08 pketa = -1.110223025e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.792752505e-01 lpclm = -1.048758818e-8
+ pdiblc1 = 5.315421921e-01 lpdiblc1 = -3.163481747e-8
+ pdiblc2 = 2.737215973e-02 lpdiblc2 = -4.685097180e-09 ppdiblc2 = -2.775557562e-29
+ pdiblcb = 1.891439592e+00 lpdiblcb = -5.432629582e-07 wpdiblcb = -7.105427358e-21
+ drout = -6.783326782e-01 ldrout = 3.008663122e-7
+ pscbe1 = 7.999049073e+08 lpscbe1 = 1.704680709e-2
+ pscbe2 = 1.829494379e-08 lpscbe2 = -2.355610367e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.033382372e+01 lbeta0 = -3.549228047e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.647441449e-09 lagidl = 6.601932258e-16 wagidl = -6.436499141e-30 pagidl = -4.846761402e-37
+ bgidl = 1.854155600e+09 lbgidl = -1.531201959e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.593976841e-01 lkt1 = -4.074556472e-8
+ kt2 = -5.800457968e-02 lkt2 = 1.294032692e-9
+ at = 1.949294486e+05 lat = -3.166706240e-2
+ ute = -1.734341181e+00 lute = 2.242768531e-7
+ ua1 = 1.543285759e-10 lua1 = 3.507348664e-17
+ ub1 = -3.113283727e-19 lub1 = 3.539735529e-26
+ uc1 = -2.735273461e-10 luc1 = 4.378123603e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.161 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {7.309927222e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.648500067e-06 wvth0 = -5.596593267e-06 pvth0 = 1.098415378e-12
+ k1 = 3.173512274e-01 lk1 = 1.480519562e-07 wk1 = 5.026303899e-07 pk1 = -9.864875346e-14
+ k2 = -2.097217495e+00 lk2 = 3.702762832e-07 wk2 = 1.257073450e-06 pk2 = -2.467195207e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.803382218e+00 ldsub = 1.027911341e-06 wdsub = 3.489718681e-06 pdsub = -6.849096369e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {2.583017024e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.141606183e-06 wvoff = -1.745555194e-05 pvoff = 3.425913901e-12
+ nfactor = {-3.846640418e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.614349572e-05 wnfactor = 2.585041911e-04 pnfactor = -5.073532507e-11
+ eta0 = -1.021668536e+01 leta0 = 2.101347602e-06 weta0 = 7.133992937e-06 peta0 = -1.400153124e-12
+ etab = -6.088076025e-01 letab = 1.193204603e-07 wetab = 4.050882592e-07 petab = -7.950464719e-14
+ u0 = -2.588277479e-01 lu0 = 5.142434751e-08 wu0 = 1.745836388e-07 pu0 = -3.426465787e-14
+ ua = -2.528058214e-08 lua = 4.511649890e-15 wua = 1.531687442e-14 pua = -3.006166358e-21
+ ub = -2.706933495e-17 lub = 5.729712475e-24 wub = 1.945215094e-23 pub = -3.817776405e-30
+ uc = 4.556542209e-10 luc = -9.204565946e-17 wuc = -3.124914091e-16 puc = 6.133112641e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.138674478e+06 lvsat = -2.100945145e-01 wvsat = -7.132626604e-01 pvsat = 1.399884960e-7
+ a0 = 5.656738450e+00 la0 = -9.380698116e-07 wa0 = -3.184709559e-06 pa0 = 6.250470215e-13
+ ags = 1.250000060e+00 lags = -1.009269113e-14 wags = -2.619970019e-15 pags = 5.142055670e-22
+ a1 = 0.0
+ a2 = 8.055819767e+00 la2 = -1.434133067e-06 wa2 = -4.868825648e-06 pa2 = 9.555800659e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.869858104e+00 lketa = -3.694520033e-07 wketa = -1.254275090e-06 pketa = 2.461703004e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.606457327e-01 lpclm = -7.825821410e-09 wpclm = -2.656834501e-08 ppclm = 5.214436233e-15
+ pdiblc1 = -6.075781447e+00 lpdiblc1 = 1.262151574e-06 wpdiblc1 = 4.284955466e-06 ppdiblc1 = -8.409867845e-13
+ pdiblc2 = 3.216798682e-02 lpdiblc2 = -6.070645791e-09 wpdiblc2 = -2.060960910e-08 ppdiblc2 = 4.044944930e-15
+ pdiblcb = 3.623729204e+01 lpdiblcb = -7.335670224e-06 wpdiblcb = -2.490431356e-05 ppdiblcb = 4.887845101e-12
+ drout = 1.000000040e+00 ldrout = -2.856694437e-15 wdrout = 8.593150369e-14 pdrout = -1.686535001e-20
+ pscbe1 = 1.240636410e+08 lpscbe1 = 1.326626495e+02 wpscbe1 = 4.503845075e+02 ppscbe1 = -8.839471537e-5
+ pscbe2 = 1.467024817e-07 lpscbe2 = -2.778090227e-14 wpscbe2 = -9.431507914e-14 ppscbe2 = 1.851074901e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -4.345903766e+00 lbeta0 = 2.492535986e-06 wbeta0 = 8.462061670e-06 pbeta0 = -1.660806534e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.755571606e-07 lagidl = 7.391192649e-14 wagidl = 2.509280990e-13 pagidl = -4.924840335e-20
+ bgidl = 1.000000386e+09 lbgidl = -6.710067749e-05 wbgidl = -6.667907715e-05 pbgidl = 1.308676910e-11
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.876691714e-02 lkt1 = -9.968753231e-08 wkt1 = -3.384354329e-07 pkt1 = 6.642303023e-14
+ kt2 = -1.539395024e+00 lkt2 = 2.921618435e-07 wkt2 = 9.918779102e-07 pkt2 = -1.946709180e-13
+ at = 1.334630430e+06 lat = -2.583535160e-01 wat = -8.771000634e-01 pat = 1.721440439e-7
+ ute = 1.075885496e+01 lute = -2.206431738e-06 wute = -7.490749621e-06 pute = 1.470171974e-12
+ ua1 = 1.417560805e-08 lua1 = -2.713486851e-15 wua1 = -9.212181046e-15 pua1 = 1.808028713e-21
+ ub1 = -1.885469845e-17 lub1 = 3.678168674e-24 wub1 = 1.248723840e-23 pub1 = -2.450807845e-30
+ uc1 = -4.540808258e-10 luc1 = 8.336941261e-17 wuc1 = 2.830358976e-16 puc1 = -5.555004044e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.162 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.163 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.120472155e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.870888723e-7
+ k1 = 4.170862753e-01 lk1 = 2.913759846e-7
+ k2 = 2.448249051e-02 lk2 = -5.836714509e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = -4.235164736e-28 pcit = 5.082197684e-32
+ voff = {-2.688785328e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.293878253e-7
+ nfactor = {2.183144685e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.000922662e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.113674562e-02 lu0 = -1.256245066e-8
+ ua = -9.216113352e-10 lua = 2.090566673e-15
+ ub = 1.520604476e-18 lub = -5.620003986e-24
+ uc = -1.046565291e-10 luc = -2.012847738e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.288282795e+04 lvsat = -2.545272048e-1
+ a0 = 1.626037978e+00 la0 = -3.240640463e-6
+ ags = 1.127453634e-01 lags = 1.089233216e-8
+ a1 = 0.0
+ a2 = 1.083322921e+00 la2 = -2.266375124e-06 wa2 = 8.881784197e-22
+ b0 = -2.350169889e-07 lb0 = 2.106462362e-12
+ b1 = 4.206262362e-10 lb1 = 3.533945400e-15
+ keta = 3.418087999e-02 lketa = -2.163844674e-07 wketa = 2.775557562e-23
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.896493835e-02 lpclm = 1.679237053e-06 wpclm = -1.387778781e-23 ppclm = 1.110223025e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.907724688e-03 lpdiblc2 = -1.261085430e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.864397580e-09 lpscbe2 = 2.392366917e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.666054167e-11 lalpha0 = 1.333161838e-15
+ alpha1 = -6.666054167e-11 lalpha1 = 1.333161838e-15
+ beta0 = 4.799834625e+01 lbeta0 = -3.599536962e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.809193870e-09 lagidl = -1.817806134e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443729441e-01 lkt1 = 1.224543810e-7
+ kt2 = -6.520326764e-02 lkt2 = 1.331404597e-07 wkt2 = 5.551115123e-23
+ at = 7.714160610e+04 lat = -1.230276006e-1
+ ute = 5.604140827e-01 lute = -1.286740876e-05 wute = 1.110223025e-22 pute = 8.881784197e-28
+ ua1 = 3.770448273e-09 lua1 = -3.360373048e-14 wua1 = 3.308722450e-30
+ ub1 = -2.644626951e-18 lub1 = 2.831349847e-23
+ uc1 = -9.425493132e-11 luc1 = 1.289271244e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.164 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.074934676e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.282250820e-8
+ k1 = 4.603687398e-01 lk1 = -5.485191820e-8
+ k2 = 1.663300362e-02 lk2 = 4.422980655e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.526831662e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.983679658e-8
+ nfactor = {1.083406992e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.796170572e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.366897430e-03 lu0 = 9.594299004e-9
+ ua = -8.793373383e-10 lua = 1.752405770e-15
+ ub = 9.308044156e-19 lub = -9.020370027e-25
+ uc = -1.070081003e-10 luc = -1.317636749e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.342668478e+04 lvsat = -1.889970965e-2
+ a0 = 1.169514648e+00 la0 = 4.112106358e-7
+ ags = 4.518586659e-02 lags = 5.513186502e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.904470373e-08 lb0 = 7.415555649e-14
+ b1 = 2.692493660e-09 lb1 = -1.463932417e-14 pb1 = -6.617444900e-36
+ keta = 7.537928491e-03 lketa = -3.260437949e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.076066625e-01 lpclm = 4.388121945e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.324642703e-04 lpdiblc2 = 7.899977302e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.461814170e-08 lpscbe2 = -2.210205481e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.999816250e-10 lalpha0 = -7.997795135e-16
+ alpha1 = 1.999816250e-10 lalpha1 = -7.997795135e-16
+ beta0 = -2.399503875e+01 lbeta0 = 2.159404686e-04 wbeta0 = -3.552713679e-21 pbeta0 = 4.263256415e-26
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.936827142e-10 lagidl = -1.255526991e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.138822703e-01 lkt1 = -1.214485986e-7
+ kt2 = -3.857419708e-02 lkt2 = -7.987253241e-8
+ at = 2.254069419e+04 lat = 3.137395630e-1
+ ute = -1.913180623e+00 lute = 6.919530795e-6
+ ua1 = -2.950544819e-09 lua1 = 2.015927433e-14
+ ub1 = 2.918299229e-18 lub1 = -1.618582223e-23 wub1 = 1.540743956e-39 pub1 = 6.162975822e-45
+ uc1 = 5.518884344e-10 luc1 = -3.879400767e-15 puc1 = -1.654361225e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.165 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.073354483e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.650289888e-8
+ k1 = 3.860761503e-01 lk1 = 2.422638348e-7
+ k2 = 3.864608706e-02 lk2 = -8.361317351e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.598897400e-01 ldsub = -1.199338541e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.344875018e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.706751263e-8
+ nfactor = {2.301599641e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.570464991e-8
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394744587e-01 letab = 2.778467713e-7
+ u0 = 1.198857651e-02 lu0 = -4.889755366e-9
+ ua = -1.319018025e-10 lua = -1.236787009e-15
+ ub = 5.490351914e-19 lub = 6.247592937e-25
+ uc = -1.334915649e-10 luc = 1.045967563e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.358762876e+04 lvsat = -9.952866729e-2
+ a0 = 1.399225751e+00 la0 = -5.074649400e-7
+ ags = -4.159569572e-02 lags = 8.983811150e-07 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.819412950e-08 lb0 = 7.755722824e-14
+ b1 = -2.575139163e-09 lb1 = 6.427335412e-15
+ keta = 2.261809468e-02 lketa = -6.357001880e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.069927487e-01 lpclm = 3.304700303e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.186804914e-04 lpdiblc2 = 4.526971437e-11
+ pdiblcb = -4.249265000e-01 lpdiblcb = 7.995590540e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.717023012e-09 lpscbe2 = 1.498082628e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.996325000e-11 lalpha0 = 3.997795270e-16
+ alpha1 = -9.996325000e-11 lalpha1 = 3.997795270e-16
+ beta0 = 5.442312590e+01 lbeta0 = -9.767455261e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.805953197e-11 lagidl = 1.790882113e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.356331678e-01 lkt1 = -3.446099523e-8
+ kt2 = -6.315530546e-02 lkt2 = 1.843383399e-8
+ at = 1.619156016e+05 lat = -2.436576261e-1
+ ute = -9.264321097e-02 lute = -3.612807586e-7
+ ua1 = 2.877410594e-09 lua1 = -3.148263775e-15
+ ub1 = -1.895518164e-18 lub1 = 3.065909193e-24
+ uc1 = -8.716392777e-10 luc1 = 1.813663789e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.166 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.086028606e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.184182979e-8
+ k1 = 5.064839054e-01 lk1 = 1.536824197e-9
+ k2 = -2.175514322e-03 lk2 = -1.999974616e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000200e-01 ldsub = -1.997795529e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.136546851e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.458280866e-8
+ nfactor = {2.242862352e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.172675677e-8
+ eta0 = -4.886402175e-01 leta0 = 9.779209169e-07 weta0 = 1.856154119e-22 peta0 = -1.040834086e-28
+ etab = 2.464242746e-04 letab = -1.492299927e-9
+ u0 = 1.041902600e-02 lu0 = -1.751807974e-9
+ ua = -6.756220924e-10 lua = -1.497460633e-16
+ ub = 8.575638770e-19 lub = 7.928691116e-27
+ uc = -1.187352451e-10 luc = 7.509496275e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.581072052e+04 lvsat = 3.597533316e-2
+ a0 = 1.033650996e+00 la0 = 2.234158726e-7
+ ags = 2.513648550e-01 lags = 3.126753396e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 8.083645775e-08 lb0 = -4.768138616e-14
+ b1 = 4.795263422e-09 lb1 = -8.308052512e-15 wb1 = 1.654361225e-30 pb1 = 1.654361225e-36
+ keta = -1.731434613e-02 lketa = 1.626551248e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.164189562e-01 lpclm = -2.881549565e-07 wpclm = 8.881784197e-22
+ pdiblc1 = 3.956566993e-01 lpdiblc1 = -1.130924086e-8
+ pdiblc2 = 4.526390171e-04 lpdiblc2 = -2.262237742e-11
+ pdiblcb = 1.748530000e-01 lpdiblcb = -3.995591080e-07 wpdiblcb = 5.551115123e-23 ppdiblcb = 8.326672685e-29
+ drout = 3.837641586e-01 ldrout = 3.523421494e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.762341479e-09 lpscbe2 = -5.917859960e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.665153203e+00 lbeta0 = 1.804820678e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.216142405e-10 lagidl = 8.118944782e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.266945131e-01 lkt1 = -5.233173475e-8
+ kt2 = -5.930686777e-02 lkt2 = 1.073978722e-8
+ at = 2.833087101e+04 lat = 2.341365030e-2
+ ute = 5.008903148e-01 lute = -1.547911563e-06 pute = 4.440892099e-28
+ ua1 = 3.034530159e-09 lua1 = -3.462387422e-15 pua1 = 1.654361225e-36
+ ub1 = -1.577991139e-18 lub1 = 2.431088525e-24 pub1 = 3.851859889e-46
+ uc1 = 4.156291695e-12 luc1 = 6.271635987e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.167 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.066457169e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.228477766e-8
+ k1 = 5.809893998e-01 lk1 = -7.291390867e-8
+ k2 = -3.726522465e-02 lk2 = 3.306394477e-08 wk2 = 6.938893904e-24 pk2 = 3.469446952e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.789122000e-01 ldsub = 7.383690995e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.182236678e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.001718417e-8
+ nfactor = {1.200359609e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.083463260e-6
+ eta0 = 9.711211764e-01 leta0 = -4.807675523e-7
+ etab = -1.493584618e-03 letab = 2.464300584e-10
+ u0 = 4.964807659e-03 lu0 = 3.698401517e-9
+ ua = -1.109598808e-09 lua = 2.839116794e-16
+ ub = 2.494279967e-19 lub = 6.156175915e-25
+ uc = -3.884456477e-11 luc = -4.736997978e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.035589602e+04 lvsat = 1.144819836e-2
+ a0 = 1.399952291e+00 la0 = -1.426161911e-7
+ ags = -1.204516172e-01 lags = 6.842185266e-7
+ a1 = 0.0
+ a2 = 1.107391439e+00 la2 = -3.071655067e-07 wa2 = 8.881784197e-22
+ b0 = 6.619131360e-08 lb0 = -3.304700618e-14
+ b1 = -7.032627217e-09 lb1 = 3.511144627e-15
+ keta = 4.139479423e-02 lketa = -4.240047666e-08 wketa = 6.938893904e-24 pketa = -8.673617380e-30
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.233102479e-01 lpclm = -1.951146831e-7
+ pdiblc1 = 6.983437078e-01 lpdiblc1 = -3.137737744e-7
+ pdiblc2 = 5.691890659e-05 lpdiblc2 = 3.728068788e-10
+ pdiblcb = -0.225
+ drout = 9.604260361e-01 ldrout = -2.238958816e-07 wdrout = -8.881784197e-22
+ pscbe1 = 1.460742549e+09 lpscbe1 = -6.602569028e+02 ppscbe1 = 4.768371582e-19
+ pscbe2 = -5.973317864e-08 lpscbe2 = 6.885265491e-14 wpscbe2 = -1.323488980e-29 ppscbe2 = 1.323488980e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.503379304e+00 lbeta0 = 1.966475673e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.554343458e-09 lagidl = -3.200021832e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.742565584e-01 lkt1 = -4.804647554e-9
+ kt2 = -3.759050968e-02 lkt2 = -1.096060934e-8
+ at = 2.356499624e+04 lat = 2.817602215e-2
+ ute = -1.856529547e+00 lute = 8.077755953e-7
+ ua1 = -2.523326854e-09 lua1 = 2.091384566e-15 wua1 = 8.271806126e-31 pua1 = 4.135903063e-37
+ ub1 = 2.573680751e-18 lub1 = -1.717531887e-24 wub1 = -1.540743956e-39
+ uc1 = 2.009891904e-10 luc1 = -1.339718666e-16 wuc1 = -1.033975766e-31 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.168 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.007966096e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.917767921e-9
+ k1 = 2.924500733e-01 lk1 = 7.114367819e-8
+ k2 = 7.415324063e-02 lk2 = -2.256339530e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.214775846e+00 ldsub = -1.072300629e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.351612806e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.560826904e-9
+ nfactor = {4.072480519e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.504861863e-7
+ eta0 = -4.722423533e-01 leta0 = 2.398533403e-07 weta0 = 8.326672685e-23 peta0 = 6.245004514e-29
+ etab = -1.925464442e-03 letab = 4.620525390e-10
+ u0 = 1.787885262e-02 lu0 = -2.749129141e-09 wu0 = -1.387778781e-23
+ ua = 2.200897025e-10 lua = -3.799552548e-16
+ ub = 1.376476647e-18 lub = 5.292164706e-26
+ uc = -9.553602869e-11 luc = 2.356706576e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.819169822e+04 lvsat = 1.752135658e-2
+ a0 = 1.611671360e+00 la0 = -2.483201119e-7
+ ags = 9.950076830e-01 lags = 1.273087391e-7
+ a1 = 0.0
+ a2 = 1.891834845e-01 la2 = 1.512635879e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.534929780e-02 lketa = 5.900462451e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.284134026e-01 lpclm = 1.018964903e-7
+ pdiblc1 = -2.639010008e-01 lpdiblc1 = 1.666413300e-07 wpdiblc1 = -1.110223025e-22 ppdiblc1 = -2.775557562e-29
+ pdiblc2 = -6.946398880e-03 lpdiblc2 = 3.869318333e-09 wpdiblc2 = 2.602085214e-24 ppdiblc2 = 1.301042607e-30
+ pdiblcb = -1.621654265e-01 lpdiblcb = -3.137110336e-8
+ drout = 4.953180247e-01 ldrout = 8.316269749e-9
+ pscbe1 = -5.214584712e+08 lpscbe1 = 3.293866893e+02 ppscbe1 = 1.192092896e-19
+ pscbe2 = 1.473011627e-07 lpscbe2 = -3.451234553e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.975670309e+00 lbeta0 = 2.328823045e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.822993481e-09 lagidl = -4.541297369e-16
+ bgidl = 7.608364006e+08 lbgidl = 1.194060145e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.450140790e-01 lkt1 = -1.940439406e-8
+ kt2 = -6.625502520e-02 lkt2 = 3.350579994e-9
+ at = 9.207669362e+04 lat = -6.029470441e-3
+ ute = 3.556362895e-01 lute = -2.966813811e-7
+ ua1 = 3.032134340e-09 lua1 = -6.822627670e-16
+ ub1 = -1.561509020e-18 lub1 = 3.470236344e-25
+ uc1 = -3.690176234e-11 luc1 = -1.520124011e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.169 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.981652160e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.428728428e-8
+ k1 = -6.868110801e-01 lk1 = 3.152392096e-7
+ k2 = 4.810608589e-01 lk2 = -1.239912228e-07 wk2 = -1.665334537e-22 pk2 = 1.387778781e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.682474392e+00 ldsub = -2.238109408e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {8.041300560e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.022245136e-8
+ nfactor = {1.047285534e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.035890417e-7
+ eta0 = 4.900000008e-01 leta0 = -5.696021432e-17
+ etab = 1.925516612e-03 letab = -4.978622536e-10 wetab = -6.505213035e-25
+ u0 = 1.623006395e-02 lu0 = -2.338143833e-9
+ ua = 1.228104028e-09 lua = -6.312179456e-16
+ ub = 2.170685950e-19 lub = 3.419214952e-25
+ uc = 3.061872191e-11 luc = -7.878898151e-18 wuc = 3.231174268e-33 puc = 8.077935669e-40
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.760102185e+05 lvsat = -1.932462687e-2
+ a0 = -5.465138832e-02 la0 = 1.670358279e-7
+ ags = 2.160686824e+00 lags = -1.632542721e-7
+ a1 = 0.0
+ a2 = 9.172257814e-01 la2 = -3.021187522e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.064756593e-02 lketa = 1.220643526e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.792752505e-01 lpclm = -1.048758818e-8
+ pdiblc1 = 5.315421921e-01 lpdiblc1 = -3.163481747e-8
+ pdiblc2 = 2.737215973e-02 lpdiblc2 = -4.685097180e-9
+ pdiblcb = 1.891439592e+00 lpdiblcb = -5.432629582e-07 wpdiblcb = -8.881784197e-22
+ drout = -6.783326782e-01 ldrout = 3.008663122e-7
+ pscbe1 = 7.999049073e+08 lpscbe1 = 1.704680709e-2
+ pscbe2 = 1.829494379e-08 lpscbe2 = -2.355610367e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.033382372e+01 lbeta0 = -3.549228047e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.647441449e-09 lagidl = 6.601932258e-16 wagidl = -6.914712933e-31 pagidl = 1.361132160e-37
+ bgidl = 1.854155600e+09 lbgidl = -1.531201959e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.593976841e-01 lkt1 = -4.074556472e-8
+ kt2 = -5.800457968e-02 lkt2 = 1.294032692e-9
+ at = 1.949294486e+05 lat = -3.166706240e-2
+ ute = -1.734341181e+00 lute = 2.242768531e-7
+ ua1 = 1.543285759e-10 lua1 = 3.507348664e-17
+ ub1 = -3.113283727e-19 lub1 = 3.539735529e-26
+ uc1 = -2.735273461e-10 luc1 = 4.378123603e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.170 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-2.035540184e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.856880933e-07 wvth0 = 5.369491373e-07 pvth0 = -1.053843224e-13
+ k1 = 3.085815365e-01 lk1 = 1.497731396e-07 wk1 = 5.083860432e-07 pk1 = -9.977838677e-14
+ k2 = -2.324277681e-04 lk2 = -4.128849104e-08 wk2 = -1.192030133e-07 pk2 = 2.339537941e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.864269520e+00 ldsub = 1.039861387e-06 wdsub = 3.529679748e-06 pdsub = -6.927525957e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.072590444e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.309941412e-07 wvoff = 1.513676729e-06 pvoff = -2.970817632e-13
+ nfactor = {5.319763515e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.793426302e-06 wnfactor = -2.886968179e-05 pnfactor = 5.666108096e-12
+ eta0 = -1.034115755e+01 leta0 = 2.125777137e-06 weta0 = 7.215685531e-06 peta0 = -1.416186521e-12
+ etab = -6.158753654e-01 letab = 1.207076147e-07 wetab = 4.097269168e-07 petab = -8.041505332e-14
+ u0 = 6.981470448e-02 lu0 = -1.307666340e-08 wu0 = -4.110834637e-08 pu0 = 8.068129600e-15
+ ua = 1.155143520e-08 lua = -2.717185992e-15 wua = -8.856420542e-15 pua = 1.738205378e-21
+ ub = -8.318767048e-19 lub = 5.802177321e-25 wub = 2.232192246e-24 pub = -4.381012111e-31
+ uc = 4.611064477e-10 luc = -9.311574074e-17 wuc = -3.160697710e-16 puc = 6.203343360e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.742315036e+05 lvsat = 1.064624780e-01 wvsat = 3.453068903e-01 pvsat = -6.777165682e-8
+ a0 = 5.712304405e+00 la0 = -9.489754637e-07 wa0 = -3.221178162e-06 pa0 = 6.322045319e-13
+ ags = 1.250000056e+00 lags = -9.224518038e-15 wags = 2.832578616e-16 pags = -5.559375182e-23
+ a1 = 0.0
+ a2 = 8.140769462e+00 la2 = -1.450805718e-06 wa2 = -4.924579153e-06 pa2 = 9.665225274e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.891742094e+00 lketa = -3.737470646e-07 wketa = -1.268637815e-06 pketa = 2.489892007e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.611092926e-01 lpclm = -7.916801976e-09 wpclm = -2.687258487e-08 ppclm = 5.274147870e-15
+ pdiblc1 = -6.150543759e+00 lpdiblc1 = 1.276824799e-06 wpdiblc1 = 4.334022868e-06 ppdiblc1 = -8.506169982e-13
+ pdiblc2 = 3.252756969e-02 lpdiblc2 = -6.141219321e-09 wpdiblc2 = -2.084560765e-08 ppdiblc2 = 4.091263185e-15
+ pdiblcb = 3.667181665e+01 lpdiblcb = -7.420952198e-06 wpdiblcb = -2.518949728e-05 ppdiblcb = 4.943816684e-12
+ drout = 1.000000186e+00 ldrout = -3.133212978e-14 wdrout = -9.290573644e-15 pdrout = 1.823414308e-21
+ pscbe1 = 1.162055541e+08 lpscbe1 = 1.342049169e+02 wpscbe1 = 4.555418642e+02 ppscbe1 = -8.940692398e-5
+ pscbe2 = 1.483480293e-07 lpscbe2 = -2.810386567e-14 wpscbe2 = -9.539507177e-14 ppscbe2 = 1.872271376e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -4.493547100e+00 lbeta0 = 2.521513205e-06 wbeta0 = 8.558961762e-06 pbeta0 = -1.679824630e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.948766734e-08 lagidl = -9.509496672e-15 wagidl = -2.803392214e-14 pagidl = 5.502077729e-21
+ bgidl = 1.000000273e+09 lbgidl = -4.500499344e-05 wbgidl = 7.209079742e-06 pbgidl = -1.414890289e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.286210130e-02 lkt1 = -1.008464410e-07 wkt1 = -3.423108344e-07 pkt1 = 6.718363591e-14
+ kt2 = -1.556700781e+00 lkt2 = 2.955583580e-07 wkt2 = 1.003235886e-06 pkt2 = -1.969000912e-13
+ at = 1.349933649e+06 lat = -2.613570023e-01 wat = -8.871437495e-01 pat = 1.741152680e-7
+ ute = 1.088955146e+01 lute = -2.232082887e-06 wute = -7.576527302e-06 pute = 1.487007131e-12
+ ua1 = 1.433634230e-08 lua1 = -2.745033360e-15 wua1 = -9.317672866e-15 pua1 = 1.828733065e-21
+ ub1 = -1.907256693e-17 lub1 = 3.720928630e-24 wub1 = 1.263022810e-23 pub1 = -2.478871718e-30
+ uc1 = -4.590191362e-10 luc1 = 8.433863011e-17 wuc1 = 2.862769700e-16 puc1 = -5.618614951e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.171 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.172 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.120472155e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.870888723e-7
+ k1 = 4.170862753e-01 lk1 = 2.913759846e-7
+ k2 = 2.448249051e-02 lk2 = -5.836714509e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = 1.016439537e-26 pcit = -5.421010862e-32
+ voff = {-2.688785328e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.293878253e-7
+ nfactor = {2.183144685e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.000922662e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.113674562e-02 lu0 = -1.256245066e-8
+ ua = -9.216113352e-10 lua = 2.090566673e-15
+ ub = 1.520604476e-18 lub = -5.620003986e-24
+ uc = -1.046565291e-10 luc = -2.012847738e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.288282795e+04 lvsat = -2.545272048e-1
+ a0 = 1.626037978e+00 la0 = -3.240640463e-6
+ ags = 1.127453634e-01 lags = 1.089233216e-8
+ a1 = 0.0
+ a2 = 1.083322921e+00 la2 = -2.266375124e-6
+ b0 = -2.350169889e-07 lb0 = 2.106462362e-12
+ b1 = 4.206262362e-10 lb1 = 3.533945400e-15
+ keta = 3.418087999e-02 lketa = -2.163844674e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.896493835e-02 lpclm = 1.679237053e-06 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.907724688e-03 lpdiblc2 = -1.261085430e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.864397580e-09 lpscbe2 = 2.392366917e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.666054167e-11 lalpha0 = 1.333161838e-15
+ alpha1 = -6.666054167e-11 lalpha1 = 1.333161838e-15
+ beta0 = 4.799834625e+01 lbeta0 = -3.599536962e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.809193870e-09 lagidl = -1.817806134e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.443729441e-01 lkt1 = 1.224543810e-7
+ kt2 = -6.520326764e-02 lkt2 = 1.331404597e-7
+ at = 7.714160610e+04 lat = -1.230276006e-01 wat = 4.656612873e-16
+ ute = 5.604140827e-01 lute = -1.286740876e-05 wute = 1.776356839e-21 pute = 2.842170943e-26
+ ua1 = 3.770448273e-09 lua1 = -3.360373048e-14 wua1 = -1.323488980e-29
+ ub1 = -2.644626951e-18 lub1 = 2.831349847e-23 pub1 = 9.860761315e-44
+ uc1 = -9.425493132e-11 luc1 = 1.289271244e-15 wuc1 = -2.067951531e-31 puc1 = 1.654361225e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.173 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.074934676e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.282250820e-8
+ k1 = 4.603687398e-01 lk1 = -5.485191820e-8
+ k2 = 1.663300362e-02 lk2 = 4.422980655e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.526831662e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.983679658e-8
+ nfactor = {1.083406992e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.796170572e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.366897430e-03 lu0 = 9.594299004e-9
+ ua = -8.793373383e-10 lua = 1.752405770e-15
+ ub = 9.308044156e-19 lub = -9.020370027e-25 wub = -6.162975822e-39
+ uc = -1.070081003e-10 luc = -1.317636749e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.342668478e+04 lvsat = -1.889970965e-2
+ a0 = 1.169514648e+00 la0 = 4.112106358e-7
+ ags = 4.518586659e-02 lags = 5.513186502e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.904470373e-08 lb0 = 7.415555649e-14
+ b1 = 2.692493660e-09 lb1 = -1.463932417e-14
+ keta = 7.537928491e-03 lketa = -3.260437949e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.076066625e-01 lpclm = 4.388121945e-06 ppclm = -7.105427358e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 2.324642703e-04 lpdiblc2 = 7.899977302e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.461814170e-08 lpscbe2 = -2.210205481e-14 wpscbe2 = -1.058791184e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.999816250e-10 lalpha0 = -7.997795135e-16
+ alpha1 = 1.999816250e-10 lalpha1 = -7.997795135e-16
+ beta0 = -2.399503875e+01 lbeta0 = 2.159404686e-04 pbeta0 = -2.273736754e-25
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.936827142e-10 lagidl = -1.255526991e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.138822703e-01 lkt1 = -1.214485986e-7
+ kt2 = -3.857419708e-02 lkt2 = -7.987253241e-8
+ at = 2.254069419e+04 lat = 3.137395630e-1
+ ute = -1.913180623e+00 lute = 6.919530795e-6
+ ua1 = -2.950544819e-09 lua1 = 2.015927433e-14 wua1 = -3.308722450e-30 pua1 = 3.970466940e-35
+ ub1 = 2.918299229e-18 lub1 = -1.618582223e-23 pub1 = -4.930380658e-44
+ uc1 = 5.518884344e-10 luc1 = -3.879400767e-15 puc1 = 9.926167351e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.174 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.073354483e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.650289888e-8
+ k1 = 3.860761503e-01 lk1 = 2.422638348e-7
+ k2 = 3.864608706e-02 lk2 = -8.361317351e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.598897400e-01 ldsub = -1.199338541e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.344875018e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.706751263e-8
+ nfactor = {2.301599641e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.570464991e-8
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394744587e-01 letab = 2.778467713e-7
+ u0 = 1.198857651e-02 lu0 = -4.889755366e-9
+ ua = -1.319018025e-10 lua = -1.236787009e-15
+ ub = 5.490351914e-19 lub = 6.247592937e-25
+ uc = -1.334915649e-10 luc = 1.045967563e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.358762876e+04 lvsat = -9.952866729e-2
+ a0 = 1.399225751e+00 la0 = -5.074649400e-7
+ ags = -4.159569572e-02 lags = 8.983811150e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.819412950e-08 lb0 = 7.755722824e-14
+ b1 = -2.575139163e-09 lb1 = 6.427335412e-15 pb1 = -2.646977960e-35
+ keta = 2.261809468e-02 lketa = -6.357001880e-08 wketa = -5.551115123e-23
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.069927487e-01 lpclm = 3.304700303e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.186804914e-04 lpdiblc2 = 4.526971437e-11
+ pdiblcb = -4.249265000e-01 lpdiblcb = 7.995590540e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.717023012e-09 lpscbe2 = 1.498082628e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.996325000e-11 lalpha0 = 3.997795270e-16
+ alpha1 = -9.996325000e-11 lalpha1 = 3.997795270e-16
+ beta0 = 5.442312590e+01 lbeta0 = -9.767455261e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.805953197e-11 lagidl = 1.790882113e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.356331678e-01 lkt1 = -3.446099523e-8
+ kt2 = -6.315530546e-02 lkt2 = 1.843383399e-8
+ at = 1.619156016e+05 lat = -2.436576261e-1
+ ute = -9.264321098e-02 lute = -3.612807586e-7
+ ua1 = 2.877410594e-09 lua1 = -3.148263775e-15
+ ub1 = -1.895518164e-18 lub1 = 3.065909193e-24
+ uc1 = -8.716392777e-10 luc1 = 1.813663789e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.175 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.086028606e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.184182979e-8
+ k1 = 5.064839054e-01 lk1 = 1.536824197e-9
+ k2 = -2.175514322e-03 lk2 = -1.999974616e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000200e-01 ldsub = -1.997795707e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.136546851e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.458280866e-8
+ nfactor = {2.242862352e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.172675677e-8
+ eta0 = -4.886402175e-01 leta0 = 9.779209169e-07 weta0 = 7.424616477e-22 peta0 = 8.049116929e-28
+ etab = 2.464242746e-04 letab = -1.492299927e-9
+ u0 = 1.041902600e-02 lu0 = -1.751807974e-9
+ ua = -6.756220924e-10 lua = -1.497460633e-16
+ ub = 8.575638770e-19 lub = 7.928691116e-27
+ uc = -1.187352451e-10 luc = 7.509496275e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.581072052e+04 lvsat = 3.597533316e-2
+ a0 = 1.033650996e+00 la0 = 2.234158726e-7
+ ags = 2.513648550e-01 lags = 3.126753396e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 8.083645775e-08 lb0 = -4.768138616e-14
+ b1 = 4.795263422e-09 lb1 = -8.308052512e-15 wb1 = -1.323488980e-29 pb1 = -1.985233470e-35
+ keta = -1.731434613e-02 lketa = 1.626551248e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.164189562e-01 lpclm = -2.881549565e-7
+ pdiblc1 = 3.956566993e-01 lpdiblc1 = -1.130924086e-8
+ pdiblc2 = 4.526390171e-04 lpdiblc2 = -2.262237742e-11
+ pdiblcb = 1.748530000e-01 lpdiblcb = -3.995591080e-07 ppdiblcb = 6.661338148e-28
+ drout = 3.837641586e-01 ldrout = 3.523421494e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.762341479e-09 lpscbe2 = -5.917859960e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.665153203e+00 lbeta0 = 1.804820678e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.216142405e-10 lagidl = 8.118944782e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.266945131e-01 lkt1 = -5.233173475e-8
+ kt2 = -5.930686777e-02 lkt2 = 1.073978722e-8
+ at = 2.833087101e+04 lat = 2.341365030e-2
+ ute = 5.008903148e-01 lute = -1.547911563e-6
+ ua1 = 3.034530159e-09 lua1 = -3.462387422e-15
+ ub1 = -1.577991139e-18 lub1 = 2.431088525e-24 pub1 = -3.081487911e-45
+ uc1 = 4.156291695e-12 luc1 = 6.271635987e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.176 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.066457169e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.228477766e-8
+ k1 = 5.809893998e-01 lk1 = -7.291390867e-8
+ k2 = -3.726522465e-02 lk2 = 3.306394477e-08 pk2 = 5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.789122000e-01 ldsub = 7.383690995e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.182236678e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.001718417e-8
+ nfactor = {1.200359609e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.083463260e-6
+ eta0 = 9.711211764e-01 leta0 = -4.807675523e-7
+ etab = -1.493584618e-03 letab = 2.464300584e-10
+ u0 = 4.964807659e-03 lu0 = 3.698401517e-9
+ ua = -1.109598808e-09 lua = 2.839116794e-16
+ ub = 2.494279967e-19 lub = 6.156175915e-25
+ uc = -3.884456477e-11 luc = -4.736997978e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.035589602e+04 lvsat = 1.144819836e-2
+ a0 = 1.399952291e+00 la0 = -1.426161911e-7
+ ags = -1.204516172e-01 lags = 6.842185266e-7
+ a1 = 0.0
+ a2 = 1.107391439e+00 la2 = -3.071655067e-7
+ b0 = 6.619131360e-08 lb0 = -3.304700618e-14
+ b1 = -7.032627217e-09 lb1 = 3.511144627e-15
+ keta = 4.139479423e-02 lketa = -4.240047666e-08 wketa = -9.714451465e-23 pketa = -6.245004514e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.233102479e-01 lpclm = -1.951146831e-7
+ pdiblc1 = 6.983437078e-01 lpdiblc1 = -3.137737744e-7
+ pdiblc2 = 5.691890659e-05 lpdiblc2 = 3.728068788e-10
+ pdiblcb = -0.225
+ drout = 9.604260361e-01 ldrout = -2.238958816e-7
+ pscbe1 = 1.460742549e+09 lpscbe1 = -6.602569028e+02 ppscbe1 = 3.814697266e-18
+ pscbe2 = -5.973317864e-08 lpscbe2 = 6.885265491e-14 wpscbe2 = 1.058791184e-28 ppscbe2 = -1.588186776e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.503379304e+00 lbeta0 = 1.966475673e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.554343458e-09 lagidl = -3.200021832e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.742565584e-01 lkt1 = -4.804647554e-9
+ kt2 = -3.759050968e-02 lkt2 = -1.096060934e-8
+ at = 2.356499624e+04 lat = 2.817602215e-2
+ ute = -1.856529547e+00 lute = 8.077755953e-7
+ ua1 = -2.523326854e-09 lua1 = 2.091384566e-15
+ ub1 = 2.573680751e-18 lub1 = -1.717531887e-24 wub1 = -1.232595164e-38
+ uc1 = 2.009891904e-10 luc1 = -1.339718666e-16 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.177 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.007966096e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.917767921e-9
+ k1 = 2.924500733e-01 lk1 = 7.114367819e-8
+ k2 = 7.415324063e-02 lk2 = -2.256339530e-08 wk2 = -2.220446049e-22
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.214775846e+00 ldsub = -1.072300629e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.351612806e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.560826904e-9
+ nfactor = {4.072480519e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.504861863e-07 wnfactor = 2.842170943e-20
+ eta0 = -4.722423533e-01 leta0 = 2.398533403e-07 weta0 = 4.440892099e-22 peta0 = -8.326672685e-29
+ etab = -1.925464442e-03 letab = 4.620525390e-10
+ u0 = 1.787885262e-02 lu0 = -2.749129141e-09 wu0 = 1.110223025e-22
+ ua = 2.200897025e-10 lua = -3.799552548e-16
+ ub = 1.376476647e-18 lub = 5.292164706e-26
+ uc = -9.553602869e-11 luc = 2.356706576e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.819169822e+04 lvsat = 1.752135658e-2
+ a0 = 1.611671360e+00 la0 = -2.483201119e-7
+ ags = 9.950076830e-01 lags = 1.273087391e-7
+ a1 = 0.0
+ a2 = 1.891834845e-01 la2 = 1.512635879e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.534929780e-02 lketa = 5.900462451e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.284134026e-01 lpclm = 1.018964903e-7
+ pdiblc1 = -2.639010008e-01 lpdiblc1 = 1.666413300e-07 wpdiblc1 = -8.881784197e-22 ppdiblc1 = -2.220446049e-28
+ pdiblc2 = -6.946398880e-03 lpdiblc2 = 3.869318333e-09 wpdiblc2 = -6.938893904e-24 ppdiblc2 = 1.734723476e-30
+ pdiblcb = -1.621654265e-01 lpdiblcb = -3.137110336e-8
+ drout = 4.953180247e-01 ldrout = 8.316269749e-9
+ pscbe1 = -5.214584712e+08 lpscbe1 = 3.293866893e+02 ppscbe1 = -9.536743164e-19
+ pscbe2 = 1.473011627e-07 lpscbe2 = -3.451234553e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.975670309e+00 lbeta0 = 2.328823045e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.822993481e-09 lagidl = -4.541297369e-16
+ bgidl = 7.608364006e+08 lbgidl = 1.194060145e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.450140790e-01 lkt1 = -1.940439406e-8
+ kt2 = -6.625502520e-02 lkt2 = 3.350579994e-9
+ at = 9.207669362e+04 lat = -6.029470441e-3
+ ute = 3.556362895e-01 lute = -2.966813811e-07 pute = -4.440892099e-28
+ ua1 = 3.032134340e-09 lua1 = -6.822627670e-16 wua1 = -1.323488980e-29
+ ub1 = -1.561509020e-18 lub1 = 3.470236344e-25
+ uc1 = -3.690176234e-11 luc1 = -1.520124011e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.178 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-8.981652160e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.428728428e-8
+ k1 = -6.868110801e-01 lk1 = 3.152392096e-7
+ k2 = 4.810608589e-01 lk2 = -1.239912228e-07 wk2 = 6.661338148e-22 pk2 = -3.885780586e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.682474392e+00 ldsub = -2.238109408e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {8.041300560e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.022245136e-8
+ nfactor = {1.047285534e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.035890417e-7
+ eta0 = 4.900000008e-01 leta0 = -5.696065841e-17
+ etab = 1.925516612e-03 letab = -4.978622536e-10 wetab = -1.734723476e-24 petab = -1.084202172e-30
+ u0 = 1.623006395e-02 lu0 = -2.338143833e-9
+ ua = 1.228104028e-09 lua = -6.312179456e-16
+ ub = 2.170685950e-19 lub = 3.419214952e-25
+ uc = 3.061872191e-11 luc = -7.878898151e-18 wuc = 9.047287950e-32 puc = -2.584939414e-38
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.760102185e+05 lvsat = -1.932462687e-2
+ a0 = -5.465138832e-02 la0 = 1.670358279e-7
+ ags = 2.160686824e+00 lags = -1.632542721e-7
+ a1 = 0.0
+ a2 = 9.172257814e-01 la2 = -3.021187522e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.064756593e-02 lketa = 1.220643526e-08 wketa = 4.440892099e-22
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.792752505e-01 lpclm = -1.048758818e-8
+ pdiblc1 = 5.315421921e-01 lpdiblc1 = -3.163481747e-8
+ pdiblc2 = 2.737215973e-02 lpdiblc2 = -4.685097180e-09 wpdiblc2 = -1.110223025e-22
+ pdiblcb = 1.891439592e+00 lpdiblcb = -5.432629582e-7
+ drout = -6.783326782e-01 ldrout = 3.008663122e-7
+ pscbe1 = 7.999049073e+08 lpscbe1 = 1.704680709e-2
+ pscbe2 = 1.829494379e-08 lpscbe2 = -2.355610367e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.033382372e+01 lbeta0 = -3.549228047e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.647441449e-09 lagidl = 6.601932258e-16 wagidl = 4.859686099e-30 pagidl = 4.846761402e-38
+ bgidl = 1.854155600e+09 lbgidl = -1.531201959e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000693823767872944
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179005734008e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.593976841e-01 lkt1 = -4.074556472e-8
+ kt2 = -5.800457968e-02 lkt2 = 1.294032692e-9
+ at = 1.949294486e+05 lat = -3.166706240e-2
+ ute = -1.734341181e+00 lute = 2.242768531e-7
+ ua1 = 1.543285759e-10 lua1 = 3.507348664e-17
+ ub1 = -3.113283727e-19 lub1 = 3.539735529e-26
+ uc1 = -2.735273461e-10 luc1 = 4.378123603e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.179 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {6.931761337e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.574279340e-06 wvth0 = -4.631014337e-06 pvth0 = 9.089060289e-13
+ k1 = -2.628487722e-01 lk1 = 2.619249091e-07 wk1 = 8.377081873e-07 pk1 = -1.644127974e-13
+ k2 = -2.425176646e+00 lk2 = 4.346431860e-07 wk2 = 1.278321439e-06 pk2 = -2.508897572e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.014667199e+00 ldsub = -8.990281283e-07 wdsub = -2.163670031e-06 pdsub = 4.246526986e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.744966090e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.496805518e-06 wvoff = -1.031354298e-05 pvoff = 2.024187514e-12
+ nfactor = {-2.972626325e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.898965814e-05 wnfactor = 1.731047760e-04 pnfactor = -3.397440886e-11
+ eta0 = 7.844185518e+00 leta0 = -1.443369221e-06 weta0 = -3.264745905e-06 peta0 = 6.407553550e-13
+ etab = 4.209530705e-01 letab = -8.278551823e-08 wetab = -1.878097527e-07 petab = 3.686048112e-14
+ u0 = -3.174576055e-01 lu0 = 6.293133651e-08 wu0 = 1.820813331e-07 pu0 = -3.573619285e-14
+ ua = -5.558087809e-08 lua = 1.045853748e-14 wua = 2.983273720e-14 pua = -5.855122166e-21
+ ub = 1.046221058e-17 lub = -1.636416309e-24 wub = -4.276725786e-24 pub = 8.393715865e-31
+ uc = -4.437969043e-10 luc = 8.448511563e-17 wuc = 2.054368896e-16 puc = -4.032007114e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.603018575e+06 lvsat = -1.282554009e+00 wvsat = -3.733397257e+00 pvsat = 7.327352126e-7
+ a0 = -2.980522216e-02 la0 = 1.779996822e-07 wa0 = 8.806852152e-08 pa0 = -1.728476838e-14
+ ags = 1.249999925e+00 lags = 1.645167913e-14 wags = 7.567882676e-14 pags = -1.485310719e-20
+ a1 = 0.0
+ a2 = -6.399707107e+00 la2 = 1.402980915e-06 wa2 = 3.455271980e-06 pa2 = -6.781489551e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.392541835e+00 lketa = 2.708429208e-07 wketa = 6.241344251e-07 pketa = -1.224957429e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.639954845e-01 lpclm = -8.483260441e-09 wpclm = -2.853593193e-08 ppclm = 5.600604681e-15
+ pdiblc1 = 1.207146761e+00 lpdiblc1 = -1.672323309e-07 wpdiblc1 = 9.369752912e-08 ppdiblc1 = -1.838954555e-14
+ pdiblc2 = 2.587249478e-02 lpdiblc2 = -4.835061045e-09 wpdiblc2 = -1.701020812e-08 ppdiblc2 = 3.338508496e-15
+ pdiblcb = -1.505112984e+01 lpdiblcb = 2.730451897e-06 wpdiblcb = 4.619057460e-06 ppdiblcb = -9.065593124e-13
+ drout = 1.000000035e+00 ldrout = -1.849869591e-15 wdrout = 7.728107221e-14 pdrout = -1.516756498e-20
+ pscbe1 = 1.264277769e+09 lpscbe1 = -9.112147628e+01 wpscbe1 = -2.061059300e+02 ppscbe1 = 4.045138035e-5
+ pscbe2 = -1.183689912e-08 lpscbe2 = 3.334829308e-15 wpscbe2 = -3.078575292e-15 ppscbe2 = 6.042165797e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.759763187e+01 lbeta0 = -1.814212035e-06 wbeta0 = -4.172449771e-06 pbeta0 = 8.189058543e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.349412312e-07 lagidl = 6.594044110e-14 wagidl = 1.935170652e-13 pagidl = -3.798062681e-20
+ bgidl = 1.000000377e+09 lbgidl = -6.539665985e-05 wbgidl = -5.266894531e-05 pbgidl = 1.033706665e-11
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.641009685e-01 lkt1 = -1.669804979e-07 wkt1 = -5.365066951e-07 pkt1 = 1.052974865e-13
+ kt2 = 1.009043618e+00 lkt2 = -2.080074665e-07 wkt2 = -4.754333997e-07 pkt2 = 9.331093620e-14
+ at = -5.351897721e+05 lat = 1.086267459e-01 wat = 1.992754993e-01 pat = -3.911080588e-8
+ ute = -2.257020594e+00 lute = 3.481290776e-07 wute = -6.859134771e-14 pute = 1.346208123e-20
+ ua1 = 3.100399619e-11 lua1 = 6.260386273e-17 wua1 = -1.073334737e-15 pua1 = 2.106580421e-22
+ ub1 = 3.175901866e-18 lub1 = -6.456670971e-25 wub1 = -1.918314488e-25 pub1 = 3.764979929e-32
+ uc1 = -7.316125429e-10 luc1 = 1.378391751e-16 wuc1 = 4.433758214e-16 puc1 = -8.701915558e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.180 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.181 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.144201227e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.616528667e-07 wvth0 = 1.343805809e-08 pvth0 = -2.687512848e-13
+ k1 = 3.624829117e-01 lk1 = 1.383403124e-06 wk1 = 3.092254007e-08 pk1 = -6.184280733e-13
+ k2 = 3.970286527e-02 lk2 = -3.627634533e-07 wk2 = -8.619480871e-09 pk2 = 1.723832821e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = -4.235164736e-28 pcit = -1.355252716e-32
+ voff = {-2.819221662e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.902509070e-07 wvoff = 7.386766139e-09 pvoff = -1.477298935e-13
+ nfactor = {2.408812771e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.514118505e-06 wnfactor = -1.277985448e-07 pnfactor = 2.555876964e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.131229127e-02 lu0 = -1.607323472e-08 wu0 = -9.941361068e-11 pu0 = 1.988199145e-15
+ ua = -8.459282372e-10 lua = 5.769603393e-16 wua = -4.286024663e-17 pua = 8.571734302e-22
+ ub = 1.227742260e-18 lub = 2.370250925e-25 wub = 1.658513876e-25 pub = -3.316905852e-30
+ uc = -1.114369971e-10 luc = 1.154758980e-16 wuc = 3.839860365e-18 puc = -7.679438501e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.402172949e+05 lvsat = -1.201181753e+00 wvsat = -2.680607665e-02 pvsat = 5.361018306e-7
+ a0 = 2.060605020e+00 la0 = -1.193166190e-05 wa0 = -2.461005309e-07 pa0 = 4.921829734e-12
+ ags = 1.414132419e-01 lags = -5.624441667e-07 wags = -1.623496360e-08 pags = 3.246873394e-13
+ a1 = 0.0
+ a2 = 1.504801083e+00 la2 = -1.069562858e-05 wa2 = -2.386881409e-07 pa2 = 4.773587382e-12
+ b0 = -2.809662902e-07 lb0 = 3.025414615e-12 wb0 = 2.602164072e-14 pb0 = -5.204136884e-19
+ b1 = -4.332680511e-09 lb1 = 9.859658666e-14 wb1 = 2.691854651e-15 pb1 = -5.383511450e-20
+ keta = 7.695621445e-02 lketa = -1.071859717e-06 wketa = -2.422418521e-08 pketa = 4.844658994e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.752968433e-01 lpclm = 7.805649998e-06 wpclm = 1.734794338e-07 ppclm = -3.469461168e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 8.739304154e-03 lpdiblc2 = -1.492374224e-07 wpdiblc2 = -3.868805430e-09 ppdiblc2 = 7.737326504e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 4.530225162e+08 lpscbe1 = 6.939294647e+03 wpscbe1 = 1.964975128e+02 ppscbe1 = -3.929805830e-3
+ pscbe2 = 3.541812924e-09 lpscbe2 = 1.303714502e-13 wpscbe2 = 3.014243562e-15 ppscbe2 = -6.028265577e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.145888723e-10 lalpha0 = 6.291546223e-15 walpha0 = 1.404047888e-16 palpha0 = -2.807992578e-21
+ alpha1 = -3.145888723e-10 lalpha1 = 6.291546223e-15 walpha1 = 1.404047888e-16 palpha1 = -2.807992578e-21
+ beta0 = 1.149389955e+02 lbeta0 = -1.698717480e-03 wbeta0 = -3.790929297e-05 pbeta0 = 7.581579960e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.338288845e-09 lagidl = -2.875957195e-14 wagidl = -2.996328332e-16 pagidl = 5.992436434e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.352164212e-01 lkt1 = 3.939183653e-06 wkt1 = 1.080769512e-07 pkt1 = -2.161459587e-12
+ kt2 = -7.430426791e-02 lkt2 = 3.151537758e-07 wkt2 = 5.154005663e-09 pkt2 = -1.030763251e-13
+ at = -5.119041921e+04 lat = 2.443518582e+00 wat = 7.267596592e-02 pat = -1.453465902e-6
+ ute = 5.908096002e-01 lute = -1.347529677e-05 wute = -1.721334629e-08 pute = 3.442542740e-13
+ ua1 = 6.041680016e-09 lua1 = -7.902669599e-14 wua1 = -1.286225791e-15 pua1 = 2.572357044e-20
+ ub1 = -5.538088294e-18 lub1 = 8.618059862e-23 wub1 = 1.638601880e-24 pub1 = -3.277083322e-29
+ uc1 = -1.308907602e-10 luc1 = 2.021960895e-15 wuc1 = 2.074730955e-17 puc1 = -4.149309418e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.182 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.037731593e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.974049961e-09 wvth0 = -2.106855232e-08 pvth0 = 7.276236081e-15
+ k1 = 5.317733012e-01 lk1 = 2.920443632e-08 wk1 = -4.043726000e-08 pk1 = -4.760212224e-14
+ k2 = 2.384693164e-03 lk2 = -6.424550534e-08 wk2 = 8.068989190e-09 pk2 = 3.888778764e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.632665260e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.410194973e-07 wvoff = 5.993483643e-09 pvoff = -1.365846576e-13
+ nfactor = {-3.186986864e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.330396843e-05 wnfactor = 7.940292712e-07 pnfactor = -4.818068020e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 6.011573153e-03 lu0 = 2.632861420e-08 wu0 = 1.333848402e-09 pu0 = -9.476843510e-15
+ ua = -1.592492627e-09 lua = 6.548926734e-15 wua = 4.038683979e-16 pua = -2.716327380e-21
+ ub = 1.814382631e-18 lub = -4.455666699e-24 wub = -5.003809465e-25 pub = 2.012463141e-30
+ uc = -8.584689756e-11 luc = -8.922608957e-17 wuc = -1.198384303e-17 puc = 4.978361173e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.303759843e+04 lvsat = 6.646859513e-01 wvsat = 8.860760115e-02 pvsat = -3.871227628e-7
+ a0 = -1.821614095e-01 la0 = 6.008821102e-06 wa0 = 7.654703713e-07 pa0 = -3.169993978e-12
+ ags = -3.458985055e-03 lags = 5.964271675e-07 wags = 2.754816323e-08 pags = -2.554549467e-14
+ a1 = 0.0
+ a2 = -4.644344861e-01 la2 = 5.056808585e-06 wa2 = 7.160644227e-07 pa2 = -2.863731383e-12
+ b0 = 2.027390205e-07 lb0 = -8.438723470e-13 wb0 = -1.040282959e-13 pb0 = 5.198902181e-19
+ b1 = 3.208745678e-08 lb1 = -1.927377429e-13 wb1 = -1.664672035e-14 pb1 = 1.008592717e-19
+ keta = -9.504854437e-02 lketa = 3.040519304e-07 wketa = 5.809595062e-08 pketa = -1.740346819e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -7.773870816e-01 lpclm = 1.102207637e-05 wpclm = 2.094110887e-07 ppclm = -3.756887998e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -1.970988911e-02 lpdiblc2 = 7.833521354e-08 wpdiblc2 = 1.129359403e-08 ppdiblc2 = -4.391478626e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 1.840932451e+09 lpscbe1 = -4.162964720e+03 wpscbe1 = -5.894925384e+02 ppscbe1 = 2.357536876e-3
+ pscbe2 = 3.229640083e-08 lpscbe2 = -9.964411845e-14 wpscbe2 = -1.001141028e-14 ppscbe2 = 4.391300114e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 9.437666168e-10 lalpha0 = -3.774372799e-15 walpha0 = -4.212143663e-16 palpha0 = 1.684547873e-21
+ alpha1 = 9.437666168e-10 lalpha1 = -3.774372799e-15 walpha1 = -4.212143663e-16 palpha1 = 1.684547873e-21
+ beta0 = -2.248169865e+02 lbeta0 = 1.019080656e-03 wbeta0 = 1.137278789e-04 pbeta0 = -4.548279256e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.175722351e-09 lagidl = -2.745915948e-14 wagidl = -1.405608831e-15 pagidl = 1.483943152e-20
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.553313255e-01 lkt1 = -3.184543768e-06 wkt1 = -3.789836899e-07 pkt1 = 1.734667552e-12
+ kt2 = -1.127119628e-02 lkt2 = -1.890644679e-07 wkt2 = -1.546201699e-08 pkt2 = 6.183670337e-14
+ at = 2.959792726e+05 lat = -3.335837830e-01 wat = -1.548515482e-01 pat = 3.665869787e-7
+ ute = -1.781252181e+00 lute = 5.499454012e-06 wute = -7.471266022e-08 pute = 8.042065235e-13
+ ua1 = -9.764240049e-09 lua1 = 4.740904718e-14 wua1 = 3.858677373e-15 pua1 = -1.543187336e-20
+ ub1 = 1.159868326e-17 lub1 = -5.090097825e-23 wub1 = -4.915805639e-24 pub1 = 1.965960944e-29
+ uc1 = 2.105911446e-09 luc1 = -1.587081270e-14 wuc1 = -8.800618794e-16 puc1 = 6.790880475e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.183 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.088794810e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.141893882e-07 wvth0 = 8.744042556e-09 pvth0 = -1.119522312e-13
+ k1 = 4.392142545e-01 lk1 = 3.993725922e-07 wk1 = -3.009274610e-08 pk1 = -8.897257462e-14
+ k2 = 3.995887630e-03 lk2 = -7.068909897e-08 wk2 = 1.962282374e-08 pk2 = -7.319058498e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.598897028e-01 ldsub = -1.199338392e-06 wdsub = 2.105491292e-14 pdsub = -8.420417696e-20
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.323838213e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.175113770e-07 wvoff = -1.191339537e-09 pvoff = -1.078506457e-13
+ nfactor = {3.302472727e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.178055662e-06 wnfactor = -5.668064391e-07 pnfactor = 6.242746065e-13
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394744588e-01 letab = 2.778467713e-7
+ u0 = 1.973296072e-02 lu0 = -2.854685084e-08 wu0 = -4.385737713e-09 pu0 = 1.339729705e-14
+ ua = -9.666354216e-10 lua = 4.045957917e-15 wua = 4.727196653e-16 pua = -2.991681844e-21
+ ub = 3.987169410e-18 lub = -1.314521681e-23 wub = -1.947056665e-24 pub = 7.798102709e-30
+ uc = -9.008223656e-11 luc = -7.228784656e-17 wuc = -2.458322354e-17 puc = 1.001718732e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.753486115e+05 lvsat = -4.086616244e-01 wvsat = -5.196534563e-02 pvsat = 1.750657032e-7
+ a0 = 1.808477825e+00 la0 = -1.952272716e-06 wa0 = -2.317643606e-07 pa0 = 8.182119813e-13
+ ags = -5.920666942e-01 lags = 2.950425377e-06 wags = 3.117383321e-07 pags = -1.162097290e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -2.941835640e-07 lb0 = 1.143452753e-12 wb0 = 1.769032364e-13 pb0 = -6.036294265e-19
+ b1 = -3.377113069e-08 lb1 = 7.064820097e-14 wb1 = 1.766666436e-14 pb1 = -3.636904682e-20
+ keta = 1.277459226e-03 lketa = -8.118128439e-08 wketa = 1.208545795e-08 pketa = 9.973471040e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.673536155e+00 lpclm = -2.779080148e-06 wpclm = -1.170308329e-06 ppclm = 1.760975580e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -7.281898162e-04 lpdiblc2 = 2.422367922e-09 wpdiblc2 = 6.494864177e-10 ppdiblc2 = -1.346179240e-15
+ pdiblcb = -1.168506467e+00 lpdiblcb = 3.773332392e-06 wpdiblcb = 4.210982584e-07 ppdiblcb = -1.684083526e-12
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 4.968100619e-09 lpscbe2 = 9.648996103e-15 wpscbe2 = 2.123059739e-15 ppscbe2 = -4.615960112e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.996325000e-11 lalpha0 = 3.997795270e-16
+ alpha1 = -9.996325000e-11 lalpha1 = 3.997795270e-16
+ beta0 = 5.089053660e+01 lbeta0 = -8.354679187e-05 wbeta0 = 2.000547711e-06 pbeta0 = -8.000720440e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.001957715e-09 lagidl = 1.246285188e-15 wagidl = 2.227813748e-15 pagidl = 3.084117737e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.382172263e-01 lkt1 = 1.588773181e-06 wkt1 = 2.846193833e-07 pkt1 = -9.192569929e-13
+ kt2 = -5.681628624e-02 lkt2 = -6.917583713e-09 wkt2 = -3.589862653e-09 pkt2 = 1.435681206e-14
+ at = 2.733374498e+05 lat = -2.430331337e-01 wat = -6.309952970e-02 pat = -3.536575405e-10
+ ute = -3.485494716e+00 lute = 1.231517154e-05 wute = 1.921412522e-06 pute = -7.178827052e-12
+ ua1 = -2.717249255e-10 lua1 = 9.445963687e-15 wua1 = 1.783393234e-15 pua1 = -7.132262143e-21
+ ub1 = -1.561539222e-18 lub1 = 1.730238898e-24 wub1 = -1.891362828e-25 pub1 = 7.564061159e-31
+ uc1 = -3.698093703e-09 luc1 = 7.340941947e-15 wuc1 = 1.600655058e-15 puc1 = -3.130163948e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.184 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.035906842e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.084523253e-07 wvth0 = -2.838455631e-08 pvth0 = -3.772232294e-14
+ k1 = 6.683892763e-01 lk1 = -5.880900782e-08 wk1 = -9.168895443e-08 pk1 = 3.417456882e-14
+ k2 = -3.791164299e-02 lk2 = 1.309516024e-08 wk2 = 2.023779850e-08 pk2 = -8.548556008e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.010234519e+00 ldsub = -5.498447520e-06 wdsub = -1.557490799e-06 pdsub = 3.113836801e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.177586024e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.165481110e-08 wvoff = -5.430710237e-08 pvoff = -1.658160153e-15
+ nfactor = {4.048681120e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.669923985e-06 wnfactor = -1.022656838e-06 pnfactor = 1.535640355e-12
+ eta0 = -1.492104129e+00 leta0 = 2.984111194e-06 weta0 = 5.682736547e-07 peta0 = -1.136129628e-12
+ etab = -3.140664623e+00 letab = 6.278021224e-06 wetab = 1.778735617e-06 petab = -3.556163863e-12
+ u0 = 1.749308881e-02 lu0 = -2.406875332e-08 wu0 = -4.006126656e-09 pu0 = 1.263835395e-14
+ ua = 2.346963148e-09 lua = -2.578803728e-15 wua = -1.711726293e-15 pua = 1.375604504e-21
+ ub = -2.216318422e-18 lub = -7.428007137e-25 wub = 1.740776433e-24 pub = 4.251470707e-31
+ uc = -2.474556873e-10 luc = 2.423433855e-16 wuc = 7.289593105e-17 puc = -9.471478877e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.528290346e+05 lvsat = 2.474524571e-01 wvsat = 9.550271699e-02 pvsat = -1.197620330e-7
+ a0 = -6.729899969e-02 la0 = 1.797902237e-06 wa0 = 6.234811939e-07 pa0 = -8.916505222e-13
+ ags = 2.090936609e+00 lags = -2.413609222e-06 wags = -1.041771559e-06 pags = 1.543927663e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 3.593477169e-07 lb0 = -1.631294632e-13 wb0 = -1.577242682e-13 pb0 = 6.537963143e-20
+ b1 = 3.356741015e-08 lb1 = -6.397938688e-14 wb1 = -1.629401196e-14 pb1 = 3.152734471e-20
+ keta = -1.253380517e-01 lketa = 1.719566750e-07 wketa = 6.117512073e-08 pketa = -8.816977363e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.098038442e+00 lpclm = 3.707572864e-07 wpclm = -1.028532943e-07 ppclm = -3.731499101e-13
+ pdiblc1 = 4.116759600e-01 lpdiblc1 = -4.333598814e-08 wpdiblc1 = -9.071899576e-09 ppdiblc1 = 1.813713131e-14
+ pdiblc2 = 5.368395588e-04 lpdiblc2 = -1.067610317e-10 wpdiblc2 = -4.768377716e-11 ppdiblc2 = 4.764872958e-17
+ pdiblcb = 1.662012934e+00 lpdiblcb = -1.885625980e-06 wpdiblcb = -8.421965168e-07 ppdiblcb = 8.415775024e-13
+ drout = 7.866256700e-01 ldrout = -4.530847701e-07 wdrout = -2.281453082e-07 pdrout = 4.561229296e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.014055919e-08 lpscbe2 = -6.921192870e-16 wpscbe2 = -2.141892299e-16 ppscbe2 = 5.681994665e-23
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.412547247e-11 lalpha0 = 1.716859373e-16 walpha0 = 4.863177544e-17 palpha0 = -9.722780652e-23
+ alpha1 = -6.433066011e-10 lalpha1 = 1.486066872e-15 walpha1 = 4.209434479e-16 palpha1 = -8.415775024e-22
+ beta0 = 1.094777824e+01 lbeta0 = -3.690633067e-06 wbeta0 = -3.557925949e-06 pbeta0 = 3.112141401e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.509523112e-09 lagidl = 1.025810292e-14 wagidl = 5.057810256e-15 pagidl = -5.349501196e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.513345861e-01 lkt1 = -7.894561230e-07 wkt1 = -3.839760152e-07 pkt1 = 4.174423866e-13
+ kt2 = -8.248715580e-02 lkt2 = 4.440528732e-08 wkt2 = 1.312727527e-08 pkt2 = -1.906517669e-14
+ at = 2.071234404e+05 lat = -1.106537821e-01 wat = -1.012523775e-01 pat = 7.592399580e-8
+ ute = 6.537442114e+00 lute = -7.723335266e-06 wute = -3.418571723e-06 pute = 3.497216548e-12
+ ua1 = 8.673094252e-09 lua1 = -8.437100226e-15 wua1 = -3.193186509e-15 pua1 = 2.817239558e-21
+ ub1 = -1.117184246e-18 lub1 = 8.418555469e-25 wub1 = -2.609604733e-25 pub1 = 9.000017061e-31
+ uc1 = 3.001219790e-11 luc1 = -1.125296958e-16 wuc1 = -1.464250996e-17 puc1 = 9.924394429e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.185 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.259373095e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.436379875e-09 wvth0 = -7.957808266e-08 pvth0 = 1.343357617e-14
+ k1 = 1.025960726e+00 lk1 = -4.161176427e-07 wk1 = -2.519926018e-07 pk1 = 1.943603930e-13
+ k2 = -1.980794202e-01 lk2 = 1.731452141e-07 wk2 = 9.107100869e-08 pk2 = -7.932970379e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -8.727592563e+00 ldsub = 6.230752259e-06 wdsub = 4.671326674e-06 pdsub = -3.110402492e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.563098133e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.372206839e-08 wvoff = -1.034044294e-07 pvoff = 4.740308039e-14
+ nfactor = {-1.663586657e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.038145276e-06 wnfactor = 1.621887138e-06 pnfactor = -1.106959882e-12
+ eta0 = 4.767466953e+00 leta0 = -3.270859104e-06 weta0 = -2.149916170e-06 peta0 = 1.580062327e-12
+ etab = 6.284019093e+00 letab = -3.139735349e-06 wetab = -3.559561256e-06 petab = 1.778209361e-12
+ u0 = -3.441179329e-02 lu0 = 2.779797869e-08 wu0 = 2.229944164e-08 pu0 = -1.364787975e-14
+ ua = -2.293987935e-09 lua = 2.058736257e-15 wua = 6.707337755e-16 pua = -1.005104456e-21
+ ub = -6.281879984e-18 lub = 3.319772660e-24 wub = 3.698758085e-24 pub = -1.531395465e-30
+ uc = 1.527550966e-10 luc = -1.575732436e-16 wuc = -1.085051875e-16 puc = 8.655299990e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.528841926e+05 lvsat = -5.803607087e-02 wvsat = -6.372612468e-02 pvsat = 3.934977548e-8
+ a0 = 1.338478454e+00 la0 = 3.931580299e-07 wa0 = 3.481337156e-08 pa0 = -3.034153707e-13
+ ags = -1.896581403e+00 lags = 1.570977964e-06 wags = 1.005843611e-06 pags = -5.021825105e-13
+ a1 = 0.0
+ a2 = 2.882008062e+00 la2 = -2.080477786e-06 wa2 = -1.004986689e-06 pa2 = 1.004248024e-12
+ b0 = 3.919082662e-07 lb0 = -1.956660805e-13 wb0 = -1.844574189e-13 pb0 = 9.209313323e-20
+ b1 = -6.087329756e-08 lb1 = 3.039190691e-14 wb1 = 3.049061771e-14 pb1 = -1.522289825e-20
+ keta = 1.902207785e-01 lketa = -1.433702194e-07 wketa = -8.428194080e-08 pketa = 5.718037696e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.042421501e+00 lpclm = 4.263333487e-07 wpclm = -1.240853322e-07 ppclm = -3.519334778e-13
+ pdiblc1 = 4.552241401e-01 lpdiblc1 = -8.685216033e-08 wpdiblc1 = 1.376815286e-07 ppdiblc1 = -1.285084331e-13
+ pdiblc2 = -2.827794529e-03 lpdiblc2 = 3.255400050e-09 wpdiblc2 = 1.633647835e-09 ppdiblc2 = -1.632447104e-15
+ pdiblcb = 2.388757095e-01 lpdiblcb = -4.635347609e-07 wpdiblcb = -2.626983808e-07 ppdiblcb = 2.625052975e-13
+ drout = 1.967129753e+00 ldrout = -1.632721182e-06 wdrout = -5.701083952e-07 pdrout = 7.978346738e-13
+ pscbe1 = 3.918220285e+09 lpscbe1 = -3.115928393e+03 wpscbe1 = -1.391699132e+03 ppscbe1 = 1.390676233e-3
+ pscbe2 = -3.155295898e-07 lpscbe2 = 3.247386622e-13 wpscbe2 = 1.448605772e-13 ppscbe2 = -1.449113166e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.717490551e-10 lalpha0 = -8.574829198e-17 walpha0 = -9.726355087e-17 palpha0 = 4.856028673e-23
+ alpha1 = 1.586613202e-09 lalpha1 = -7.422139404e-16 walpha1 = -8.418868958e-16 palpha1 = 4.203246610e-22
+ beta0 = 5.043445869e+00 lbeta0 = 2.209359618e-06 wbeta0 = -3.058461765e-07 pbeta0 = -1.375480929e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.917835237e-09 lagidl = -1.160856319e-15 wagidl = -7.721617564e-16 pagidl = 4.761857875e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.677198262e-01 lkt1 = 1.289227843e-07 wkt1 = 1.095605701e-07 pkt1 = -7.573144938e-14
+ kt2 = -1.658601052e-02 lkt2 = -2.144742062e-08 wkt2 = -1.189509993e-08 pkt2 = 5.938807067e-15
+ at = 1.127524450e+05 lat = -1.635214946e-02 wat = -5.050792249e-02 pat = 2.521683792e-8
+ ute = -1.883181132e+00 lute = 6.910988217e-07 wute = 1.509311221e-08 pute = 6.607545704e-14
+ ua1 = -2.480345799e-09 lua1 = 2.708142047e-15 wua1 = -2.434068721e-17 pua1 = -3.492771626e-22
+ ub1 = 5.702864852e-19 lub1 = -8.443748932e-25 wub1 = 1.134546214e-24 pub1 = -4.944792835e-31
+ uc1 = -9.782911677e-11 luc1 = 1.521765550e-17 wuc1 = 1.692243931e-16 puc1 = -8.448781664e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.186 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-9.225465299e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.129277465e-09 wvth0 = -4.837412529e-08 pvth0 = -2.145467608e-15
+ k1 = 8.235365571e-01 lk1 = -3.150543399e-07 wk1 = -3.007606488e-07 pk1 = 2.187085720e-13
+ k2 = -1.374640911e-01 lk2 = 1.428821018e-07 wk2 = 1.198414343e-07 pk2 = -9.369377036e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.257094482e+00 ldsub = -1.250577519e-06 wdsub = -2.855525551e-06 pdsub = 6.474913846e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-6.099260215e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.930033448e-07 wvoff = 2.122337699e-07 pvoff = -1.101840252e-13
+ nfactor = {8.054465481e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.813738025e-06 wnfactor = -2.255045868e-06 pnfactor = 8.286570754e-13
+ eta0 = -4.051078263e+00 leta0 = 1.131931874e-06 weta0 = 2.026737722e-06 peta0 = -5.051947785e-13
+ etab = -9.063534744e-03 letab = 2.180549146e-09 wetab = 4.042374869e-09 petab = -9.732052503e-16
+ u0 = 2.583411440e-02 lu0 = -2.280694419e-09 wu0 = -4.505160211e-09 pu0 = -2.652802046e-16
+ ua = 2.354031079e-09 lua = -2.618569562e-16 wua = -1.208476609e-15 pua = -6.688048367e-23
+ ub = 6.950987474e-19 lub = -1.635886262e-25 wub = 3.858724812e-25 pub = 1.226123658e-31
+ uc = -3.196175834e-10 luc = 7.826590253e-17 wuc = 1.269000734e-16 puc = -3.097660765e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.472475070e+04 lvsat = 5.949452879e-03 wvsat = 1.963373984e-03 pvsat = 6.553307927e-9
+ a0 = 5.674746913e+00 la0 = -1.771789042e-06 wa0 = -2.300968443e-06 pa0 = 8.627587367e-13
+ ags = 4.662325812e-02 lags = 6.008038890e-07 wags = 5.370814804e-07 pags = -2.681459853e-13
+ a1 = 0.0
+ a2 = -4.633958195e+00 la2 = 1.671981107e-06 wa2 = 2.731403011e-06 pa2 = -8.612005797e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.491863020e-01 lketa = 2.608385661e-08 wketa = 5.314102150e-08 pketa = -1.143009831e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.854357463e+00 lpclm = -9.775678590e-07 wpclm = -2.053415633e-06 ppclm = 6.113136146e-13
+ pdiblc1 = -6.459342797e-01 lpdiblc1 = 4.629176981e-07 wpdiblc1 = 2.163500302e-07 ppdiblc1 = -1.677848626e-13
+ pdiblc2 = -8.156435988e-03 lpdiblc2 = 5.915804228e-09 wpdiblc2 = 6.852585350e-10 ppdiblc2 = -1.158949520e-15
+ pdiblcb = -8.562183106e-01 lpdiblcb = 8.320735510e-08 wpdiblcb = 3.930504769e-07 ppdiblcb = -6.488715597e-14
+ drout = -1.388758708e+00 ldrout = 4.275647016e-08 wdrout = 1.066975263e-06 pdrout = -1.950389878e-14
+ pscbe1 = -5.436431541e+09 lpscbe1 = 1.554521851e+03 wpscbe1 = 2.783408229e+03 ppscbe1 = -6.938087438e-4
+ pscbe2 = 6.617575754e-07 lpscbe2 = -1.631866144e-13 wpscbe2 = -2.913428400e-13 ppscbe2 = 7.286978253e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.067570411e+01 lbeta0 = -6.026297917e-07 wbeta0 = -1.529061541e-06 pbeta0 = 4.731605262e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.202999994e-08 lagidl = -5.710241228e-15 wagidl = -5.780350241e-15 pagidl = 2.976599011e-21
+ bgidl = -1.286768025e+08 lbgidl = 5.635088238e+02 wbgidl = 5.037420011e+02 pbgidl = -2.515007502e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.641743056e-01 lkt1 = -2.262687006e-08 wkt1 = -4.578053373e-08 pkt1 = 1.824926827e-15
+ kt2 = -2.739101506e-02 lkt2 = -1.605286003e-08 wkt2 = -2.200915531e-08 pkt2 = 1.098840092e-14
+ at = 2.298534798e+05 lat = -7.481659761e-02 wat = -7.802464735e-02 pat = 3.895497556e-8
+ ute = 1.354483266e+00 lute = -9.253536938e-07 wute = -5.656590289e-07 pute = 3.560246748e-13
+ ua1 = 5.578672842e-09 lua1 = -1.315443895e-15 wua1 = -1.442135312e-15 pua1 = 3.585780710e-22
+ ub1 = -1.239500927e-18 lub1 = 5.918861935e-26 wub1 = -1.823570471e-25 pub1 = 1.630044231e-31
+ uc1 = 1.097665386e-10 luc1 = -8.842758939e-17 wuc1 = -8.306001886e-17 puc1 = 4.146896031e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.187 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-2.859486909e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.618108378e-07 wvth0 = -3.467055647e-07 pvth0 = 7.221811864e-14
+ k1 = -6.408735257e+00 lk1 = 1.487697894e-06 wk1 = 3.240394325e-06 pk1 = -6.639774224e-13
+ k2 = 2.783241770e+00 lk2 = -5.851476445e-07 wk2 = -1.303752676e-06 pk2 = 2.611584155e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.477386114e+00 ldsub = -1.056223513e-06 wdsub = -2.149104047e-06 pdsub = 4.714052284e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.683193692e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.785911406e-07 wvoff = -9.076739362e-07 pvoff = 1.689697691e-13
+ nfactor = {-6.862920982e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.904644311e-06 wnfactor = 4.479644872e-06 pnfactor = -8.500656119e-13
+ eta0 = 4.900000036e-01 leta0 = -2.688123057e-16 weta0 = -1.607484812e-15 peta0 = 1.199741417e-22
+ etab = 9.110271781e-03 letab = -2.349544738e-09 wetab = -4.068813069e-09 petab = 1.048630011e-15
+ u0 = 6.095187998e-02 lu0 = -1.103432425e-08 wu0 = -2.532650108e-08 pu0 = 4.924751327e-15
+ ua = 1.325419297e-08 lua = -2.978885810e-15 wua = -6.810518481e-15 pua = 1.329512484e-21
+ ub = -6.434692202e-18 lub = 1.613618715e-24 wub = 3.766971960e-24 pub = -7.201773959e-31
+ uc = 1.435381904e-10 luc = -3.718262142e-17 wuc = -6.394765003e-17 puc = 1.659505013e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.144606556e+05 lvsat = -9.119806745e-02 wvsat = -1.350373439e-01 pvsat = 4.070279188e-8
+ a0 = -4.595750978e+00 la0 = 7.882866146e-07 wa0 = 2.571679191e-06 pa0 = -3.518217755e-13
+ ags = 5.547773975e+00 lags = -7.704404443e-07 wags = -1.918148098e-06 pags = 3.438568156e-13
+ a1 = 0.0
+ a2 = 2.645679952e+00 la2 = -1.425778957e-07 wa2 = -9.788443385e-07 pa2 = 6.363422578e-14
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.756443543e-01 lketa = 5.760542302e-08 wketa = 1.104290212e-07 pketa = -2.570999156e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.311145937e-01 lpclm = -4.949372529e-08 wpclm = 3.104299579e-07 ppclm = 2.208964352e-14
+ pdiblc1 = 1.810129900e+00 lpdiblc1 = -1.492931396e-07 wpdiblc1 = -7.240795620e-07 ppdiblc1 = 6.663131973e-14
+ pdiblc2 = 1.042782306e-01 lpdiblc2 = -2.211022295e-08 wpdiblc2 = -4.355283083e-08 ppdiblc2 = 9.868057825e-15
+ pdiblcb = 9.763042816e+00 lpdiblcb = -2.563802770e-06 wpdiblcb = -4.457783365e-06 ppdiblcb = 1.144255942e-12
+ drout = -6.913448850e+00 ldrout = 1.419868358e-06 wdrout = 3.531021109e-06 pdrout = -6.337042867e-13
+ pscbe1 = 7.996682030e+08 lpscbe1 = 8.044842847e-02 wpscbe1 = 1.340484605e-01 ppscbe1 = -3.590509901e-8
+ pscbe2 = 5.168451708e-08 lpscbe2 = -1.111675349e-14 wpscbe2 = -1.890891603e-14 ppscbe2 = 4.961540482e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.497773436e+01 lbeta0 = -1.674975361e-06 wbeta0 = -2.629902322e-06 pbeta0 = 7.475616035e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.337757478e-08 lagidl = 3.115627884e-15 wagidl = 1.173972327e-14 pagidl = -1.390542112e-21
+ bgidl = 5.030988053e+09 lbgidl = -7.226150364e+02 wbgidl = -1.799078340e+03 pbgidl = 3.225117621e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 3.164760679e-01 lkt1 = -1.922891854e-07 wkt1 = -3.827554163e-07 pkt1 = 8.582097092e-14
+ kt2 = -1.162913636e-01 lkt2 = 6.106885349e-09 wkt2 = 3.300850517e-08 pkt2 = -2.725576214e-15
+ at = 5.292485590e+05 lat = -1.494453120e-01 wat = -1.893289241e-01 pat = 6.669923610e-8
+ ute = -6.604018613e+00 lute = 1.058422277e-06 wute = 2.757756766e-06 pute = -4.723865633e-13
+ ua1 = -3.626547872e-10 lua1 = 1.655211364e-16 wua1 = 2.927738824e-16 pua1 = -7.387406942e-23
+ ub1 = -1.672216871e-18 lub1 = 1.670495589e-25 wub1 = 7.706874870e-25 pub1 = -7.455622274e-32
+ uc1 = -1.073885066e-09 luc1 = 2.066153278e-16 wuc1 = 4.532521811e-16 puc1 = -9.221490020e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.188 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {-1.959678017e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.513388558e-07 wvth0 = 4.043144663e-07 pvth0 = -6.833226268e-14
+ k1 = 5.054080345e+00 lk1 = -6.209707288e-07 wk1 = -2.173332575e-06 pk1 = 3.355815972e-13
+ k2 = -1.532874901e+00 lk2 = 2.064644633e-07 wk2 = 7.730002533e-07 pk2 = -1.216694084e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.400418484e-01 ldsub = 4.997042752e-09 wdsub = 9.253971595e-07 pdsub = -8.730760410e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.707365290e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.472194865e-07 wvoff = 1.101622829e-06 pvoff = -2.093611744e-13
+ nfactor = {3.275178443e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.689715238e-06 wnfactor = -1.378634850e-05 pnfactor = 2.654296432e-12
+ eta0 = 7.990146704e+00 leta0 = -1.472016292e-06 weta0 = -3.347405476e-06 peta0 = 6.569785355e-13
+ etab = 4.087775991e-01 letab = -8.101306400e-08 wetab = -1.809146372e-07 petab = 3.585671902e-14
+ u0 = 1.061984521e-02 lu0 = -2.202310888e-09 wu0 = -3.712864123e-09 pu0 = 1.149773281e-15
+ ua = -5.268156619e-09 lua = 3.739104046e-16 wua = 1.340039273e-15 pua = -1.440768399e-22
+ ub = 7.177981598e-18 lub = -9.050505450e-25 wub = -2.416827502e-24 pub = 4.251903778e-31
+ uc = -7.836650684e-10 luc = 1.412688359e-16 wuc = 3.979083093e-16 puc = -7.247737336e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.111074709e+06 lvsat = 1.995626654e-01 wvsat = 6.351863386e-01 pvsat = -1.066052453e-7
+ a0 = -7.070205820e+00 la0 = 1.348690033e-06 wa0 = 4.075131865e-06 pa0 = -6.802607625e-13
+ ags = 1.250000276e+00 lags = -4.613592619e-14 wags = -1.229633284e-13 pags = 2.059101778e-20
+ a1 = 0.0
+ a2 = 6.529191799e-01 la2 = 2.350103969e-07 wa2 = -5.387149180e-07 pa2 = -1.671323480e-14
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.039338884e+00 lketa = 2.129547487e-07 wketa = 4.241113555e-07 pketa = -8.971297642e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.344392384e+00 lpclm = 8.241980788e-07 wpclm = 2.807774218e-06 ppclm = -4.659568299e-13
+ pdiblc1 = 5.273822864e+00 lpdiblc1 = -8.432525575e-07 wpdiblc1 = -2.209309948e-06 ppdiblc1 = 3.644488210e-13
+ pdiblc2 = -1.061539971e-01 lpdiblc2 = 1.709350878e-08 wpdiblc2 = 5.775797856e-08 ppdiblc2 = -9.079903740e-15
+ pdiblcb = -3.749866367e+01 lpdiblcb = 6.468886347e-06 wpdiblcb = 1.733136524e-05 ppdiblcb = -3.023679603e-12
+ drout = 1.046127101e+00 ldrout = -7.669322852e-09 wdrout = -2.612223377e-08 pdrout = 4.343213348e-15
+ pscbe1 = 1.274257562e+09 lpscbe1 = -9.305720300e+01 wpscbe1 = -2.117576065e+02 ppscbe1 = 4.154760561e-5
+ pscbe2 = -1.129916869e-07 lpscbe2 = 2.014920135e-14 wpscbe2 = 5.420659489e-14 ppscbe2 = -8.917964079e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -9.098767740e-03 lbeta0 = 1.107574725e-06 wbeta0 = 5.798453068e-06 pbeta0 = -8.357370491e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.609257181e-08 lagidl = -1.022347023e-14 wagidl = -2.226694981e-14 pagidl = 5.151910144e-21
+ bgidl = 1.000001339e+09 lbgidl = -2.224820013e-04 wbgidl = -5.978309212e-04 pbgidl = 9.929638720e-11
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.207257862e-01 lkt1 = 1.266863118e-08 wkt1 = 7.784371408e-08 pkt1 = 3.560028924e-15
+ kt2 = 8.246197732e-01 lkt2 = -1.779819128e-07 wkt2 = -3.709919634e-07 pkt2 = 7.630710480e-14
+ at = -2.655172897e+06 lat = 4.613730159e-01 wat = 1.399847383e+00 pat = -2.388752515e-7
+ ute = -3.673634408e+00 lute = 5.836623771e-07 wute = 8.022453332e-07 pute = -1.333853205e-13
+ ua1 = 1.457407042e-09 lua1 = -1.759966520e-16 wua1 = -1.881123898e-15 pua1 = 3.457803768e-22
+ ub1 = -9.141143593e-19 lub1 = 3.410215882e-26 wub1 = 2.124393820e-24 pub1 = -3.473116876e-31
+ uc1 = -4.497806135e-11 luc1 = 2.427057194e-17 wuc1 = 5.452647485e-17 puc1 = -2.270389280e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.189 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.101117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.021564026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.25740872+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.9830912+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0105086
+ ua = -8.1707916e-10
+ ub = 1.23959395e-18
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -1.2969e-7
+ b1 = 5.97330000000002e-10
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.190 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.114092114e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.594927527e-7
+ k1 = 4.317674931e-01 lk1 = -2.237578829e-9
+ k2 = 2.039018519e-02 lk2 = 2.347595343e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.124978752e-06 lcit = 1.289879782e-10 wcit = 1.058791184e-27 pcit = 2.371692252e-32
+ voff = {-2.653714884e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.592495144e-7
+ nfactor = {2.122469260e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.787458760e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.108954662e-02 lu0 = -1.161850542e-8
+ ua = -9.419602655e-10 lua = 2.497530322e-15
+ ub = 1.599346401e-18 lub = -7.194784609e-24 wub = -7.703719778e-40
+ uc = -1.028334633e-10 luc = -5.658845390e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.509195847e+00 la0 = -9.038837261e-7
+ ags = 1.050374249e-01 lags = 1.650454355e-7
+ a1 = 0.0
+ a2 = 0.97
+ b0 = -2.226625907e-07 lb0 = 1.859383479e-12
+ b1 = 1.698648807e-09 lb1 = -2.202556667e-14 wb1 = 4.135903063e-31 pb1 = -6.617444900e-36
+ keta = 2.267986694e-02 lketa = 1.362734034e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.339858448e-02 lpclm = 3.202713342e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 7.091650036e-05 lpdiblc2 = 2.412395940e-08 ppdiblc2 = -6.938893904e-30
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.932919080e+08 lpscbe1 = -1.865769591e+3
+ pscbe2 = 1.029548202e-08 lpscbe2 = -4.696967791e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.666935995e-09 lagidl = -1.533300839e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.930608188e-01 lkt1 = -9.037504099e-7
+ kt2 = -6.275627981e-02 lkt2 = 8.420250168e-8
+ at = 1.116462644e+05 lat = -8.130954049e-1
+ ute = 5.522416336e-01 lute = -1.270396579e-05 wute = 5.551115123e-23 pute = -3.108624469e-27
+ ua1 = 3.159781723e-09 lua1 = -2.139084832e-14
+ ub1 = -1.866661400e-18 lub1 = 1.275475925e-23
+ uc1 = -8.440464839e-11 luc1 = 1.092272825e-15 wuc1 = -2.584939414e-32 puc1 = -2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.191 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.084937476e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.627707583e-8
+ k1 = 4.411701805e-01 lk1 = -7.745216767e-8
+ k2 = 2.046394981e-02 lk2 = 2.288589072e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.498376161e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.498995383e-8
+ nfactor = {1.460391437e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.508677198e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.000173957e-03 lu0 = 5.094940206e-9
+ ua = -6.875911280e-10 lua = 4.627641833e-16 wua = -4.135903063e-31
+ ub = 6.932365575e-19 lub = 5.342815071e-26
+ uc = -1.126977172e-10 luc = 2.231832719e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.054952691e+05 lvsat = -2.026955281e-1
+ a0 = 1.532940069e+00 la0 = -1.093820051e-6
+ ags = 5.826501794e-02 lags = 5.391903138e-7
+ a1 = 0.0
+ a2 = 1.139968762e+00 la2 = -1.359625173e-6
+ b0 = -3.034522532e-08 lb0 = 3.209859093e-13 wb0 = -6.617444900e-30 pb0 = 2.646977960e-35
+ b1 = -5.210936170e-09 lb1 = 3.324603460e-14 pb1 = -3.308722450e-36
+ keta = 3.512037473e-02 lketa = -8.588757816e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.081837246e-01 lpclm = 2.604449243e-06 wpclm = -4.163336342e-23 ppclm = 1.110223025e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.594368959e-03 lpdiblc2 = -2.005960053e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 5.201242759e+08 lpscbe1 = 1.119297188e+3
+ pscbe2 = 9.864984505e-09 lpscbe2 = -1.253304084e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.633620226e-11 lagidl = 5.789849111e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.938138686e-01 lkt1 = 7.021264349e-7
+ kt2 = -4.591516057e-02 lkt2 = -5.051407407e-8
+ at = -5.097879309e+04 lat = 4.877855253e-01 pat = -2.910383046e-23
+ ute = -1.948652251e+00 lute = 7.301347135e-6
+ ua1 = -1.118545169e-09 lua1 = 1.283262225e-14
+ ub1 = 5.844025759e-19 lub1 = -6.851951026e-24 pub1 = 7.703719778e-46
+ uc1 = 1.340579452e-10 luc1 = -6.552673532e-16 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.192 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.069203039e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.664910851e-8
+ k1 = 3.717888972e-01 lk1 = 2.000219706e-7
+ k2 = 4.796249337e-02 lk2 = -8.708807211e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.598897500e-01 ldsub = -1.199338581e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.350531188e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.413716868e-8
+ nfactor = {2.032494687e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.206846954e-7
+ eta0 = 1.594707838e-01 leta0 = -3.178247240e-7
+ etab = -1.394744588e-01 letab = 2.778467713e-7
+ u0 = 9.906342316e-03 lu0 = 1.470932801e-9
+ ua = 9.253319882e-11 lua = -2.657159732e-15 pua = 8.271806126e-37
+ ub = -3.753766688e-19 lub = 4.327095625e-24
+ uc = -1.451630400e-10 luc = 1.521557562e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.891583431e+04 lvsat = -1.641202499e-2
+ a0 = 1.289190061e+00 la0 = -1.189991736e-7
+ ags = 1.064095558e-01 lags = 3.466475486e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.021831847e-07 lb0 = -2.090303226e-13
+ b1 = 5.812533549e-09 lb1 = -1.083974203e-14 pb1 = -6.617444900e-36
+ keta = 2.835595576e-02 lketa = -5.883487416e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.136079455e-02 lpclm = 1.166535432e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 7.270397489e-04 lpdiblc2 = -5.938611736e-10 wpdiblc2 = -4.336808690e-25
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.724996554e-09 lpscbe2 = -6.934551689e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.996325000e-11 lalpha0 = 3.997795270e-16
+ alpha1 = -9.996325000e-11 lalpha1 = 3.997795270e-16
+ beta0 = 5.537293392e+01 lbeta0 = -1.014730866e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 9.896484883e-10 lagidl = 1.937308001e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.005032878e-01 lkt1 = -4.709003049e-7
+ kt2 = -6.485967887e-02 lkt2 = 2.525007493e-8
+ at = 1.319575862e+05 lat = -2.438255335e-1
+ ute = 8.195934769e-01 lute = -3.769601116e-06 wute = -1.110223025e-22 pute = 4.440892099e-28
+ ua1 = 3.724119314e-09 lua1 = -6.534476325e-15
+ ub1 = -1.985315152e-18 lub1 = 3.425031142e-24
+ uc1 = -1.116898904e-10 luc1 = 3.275433643e-16 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.193 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.099504855e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.393225205e-8
+ k1 = 4.629523747e-01 lk1 = 1.776202057e-8
+ k2 = 7.432866005e-03 lk2 = -6.058606654e-09 wk2 = 3.469446952e-24
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.794561000e-01 ldsub = 1.478368700e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.394382847e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.537005997e-8
+ nfactor = {1.757331485e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.708088539e-7
+ eta0 = -2.188386675e-01 leta0 = 4.385161211e-07 weta0 = -4.293440603e-23 peta0 = -2.211772432e-29
+ etab = 8.447438288e-01 letab = -1.689866403e-06 wetab = -1.791101989e-22 petab = -1.999268806e-28
+ u0 = 8.517021266e-03 lu0 = 4.248553750e-9
+ ua = -1.488305213e-09 lua = 5.033551747e-16
+ ub = 1.684039248e-18 lub = 2.097774619e-25
+ uc = -8.412615317e-11 luc = 3.012684465e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.115292645e+04 lvsat = -2.088456501e-2
+ a0 = 1.329663650e+00 la0 = -1.999166028e-7
+ ags = -2.432411841e-01 lags = 1.045692035e-6
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 5.953077744e-09 lb0 = -1.664083773e-14 wb0 = 1.654361225e-30 pb0 = 1.654361225e-36
+ b1 = -2.940709635e-09 lb1 = 6.660310706e-15 wb1 = 8.271806126e-31
+ keta = 1.173000998e-02 lketa = -2.559520267e-08 wketa = 2.602085214e-24 pketa = 5.204170428e-30
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.675868874e-01 lpclm = -4.653168279e-7
+ pdiblc1 = 3.913495973e-01 lpdiblc1 = -2.698202679e-9
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 2.754467005e-01 ldrout = 5.688974523e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.660650004e-09 lpscbe2 = -5.648093633e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.230891020e-10 lalpha0 = -4.616123357e-17
+ alpha1 = 2.998530000e-10 lalpha1 = -3.995591080e-16 walpha1 = -1.033975766e-31
+ beta0 = 2.975942507e+00 lbeta0 = 3.282384466e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.822930993e-09 lagidl = -1.727909545e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.089963376e-01 lkt1 = 1.458590524e-7
+ kt2 = -5.307437892e-02 lkt2 = 1.688137231e-9
+ at = -1.974112419e+04 lat = 5.946038866e-02 pat = 7.275957614e-24
+ ute = -1.122158620e+00 lute = 1.124758889e-7
+ ua1 = 1.518488261e-09 lua1 = -2.124835359e-15 pua1 = -4.135903063e-37
+ ub1 = -1.701888384e-18 lub1 = 2.858385925e-24 wub1 = 1.925929944e-40 pub1 = 7.703719778e-46
+ uc1 = -2.795591170e-12 luc1 = 1.098348032e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.194 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.104238773e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.866269021e-8
+ k1 = 4.613498670e-01 lk1 = 1.936335047e-8
+ k2 = 5.972921454e-03 lk2 = -4.599735162e-09 wk2 = 1.734723476e-24 pk2 = -8.673617380e-31
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.738912200e+00 ldsub = -7.383690995e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.673174013e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.248856541e-8
+ nfactor = {1.970389436e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.579075009e-7
+ eta0 = -4.960310000e-02 leta0 = 2.694049417e-7
+ etab = -1.691480682e+00 letab = 8.444939822e-7
+ u0 = 1.555200252e-02 lu0 = -2.781256795e-9
+ ua = -7.911518577e-10 lua = -1.932857728e-16
+ ub = 2.005502128e-18 lub = -1.114491425e-25
+ uc = -9.036000547e-11 luc = 3.635611507e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.010038959e+04 lvsat = 3.013044824e-2
+ a0 = 1.416480774e+00 la0 = -2.866699171e-7
+ ags = 3.570967666e-01 lags = 4.457953328e-7
+ a1 = 0.0
+ a2 = 6.302499000e-01 la2 = 1.696253337e-7
+ b0 = -2.138427100e-08 lb0 = 1.067641806e-14
+ b1 = 7.443524985e-09 lb1 = -3.716291502e-15
+ keta = 1.379920976e-03 lketa = -1.525272098e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.643977597e-01 lpclm = -3.622035443e-7
+ pdiblc1 = 7.637113163e-01 lpdiblc1 = -3.747862358e-7
+ pdiblc2 = 8.325324063e-04 lpdiblc2 = -4.022365449e-10
+ pdiblcb = -3.497223582e-01 lpdiblcb = 1.246306873e-7
+ drout = 6.897533990e-01 ldrout = 1.548952693e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.042855491e-09 lpscbe2 = 5.253107003e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.382179594e-11 lalpha0 = 2.305516105e-17
+ alpha1 = -2.997060000e-10 lalpha1 = 1.995592161e-16
+ beta0 = 4.358171495e+00 lbeta0 = 1.901171416e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.187741140e-09 lagidl = -9.392155723e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.222400495e-01 lkt1 = -4.075996989e-8
+ kt2 = -4.323799373e-02 lkt2 = -8.141018220e-9
+ at = -4.148516100e+02 lat = 4.014832089e-2
+ ute = -1.849363730e+00 lute = 8.391465037e-7
+ ua1 = -2.534883179e-09 lua1 = 1.925556854e-15 pua1 = -4.135903063e-37
+ ub1 = 3.112333783e-18 lub1 = -1.952297789e-24 wub1 = -7.703719778e-40
+ uc1 = 2.813325306e-10 luc1 = -1.740844844e-16 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.195 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.030932872e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.936380136e-9
+ k1 = 1.496567402e-01 lk1 = 1.749808194e-7
+ k2 = 1.310508365e-01 lk2 = -6.704676041e-08 wk2 = -2.081668171e-23 pk2 = 6.938893904e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.409534111e-01 ldsub = 2.001820048e-07 pdsub = -5.551115123e-29
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.343982070e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.387333611e-8
+ nfactor = {3.001843396e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.293863905e-8
+ eta0 = 0.49
+ etab = -6.25e-6
+ u0 = 1.573991974e-02 lu0 = -2.875077282e-09 wu0 = 6.938893904e-24
+ ua = -3.536635579e-10 lua = -4.117083688e-16
+ ub = 1.559678864e-18 lub = 1.111348091e-25
+ uc = -3.528717461e-11 luc = 8.860178169e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.912385712e+04 lvsat = 2.063269672e-2
+ a0 = 5.192313932e-01 la0 = 1.612952952e-7
+ ags = 1.25
+ a1 = 0.0
+ a2 = 1.485982588e+00 la2 = -2.576120468e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.011932303e-02 lketa = 4.737490779e-10
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -7.464949288e-01 lpclm = 3.921322938e-07 wpclm = 5.551115123e-23 ppclm = 7.632783294e-29
+ pdiblc1 = -1.611836339e-01 lpdiblc1 = 8.698144148e-08 wpdiblc1 = 2.775557562e-23 ppdiblc1 = -3.469446952e-30
+ pdiblc2 = -6.621055952e-03 lpdiblc2 = 3.319079247e-09 wpdiblc2 = -8.673617380e-25 ppdiblc2 = 4.336808690e-31
+ pdiblcb = 2.444471645e-02 lpdiblcb = -6.217783725e-8
+ drout = 1.001890127e+00 ldrout = -9.436740779e-10
+ pscbe1 = 8.000313575e+08 lpscbe1 = -1.565572071e-2
+ pscbe2 = 8.979160365e-09 lpscbe2 = 8.433181703e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.249711661e+00 lbeta0 = 4.575266151e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -9.213664622e-10 lagidl = 9.590820500e-16 pagidl = 2.067951531e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.667494856e-01 lkt1 = -1.853796627e-8
+ kt2 = -7.670439966e-02 lkt2 = 8.567586936e-9
+ at = 5.503262054e+04 lat = 1.246533871e-2
+ ute = 8.707609580e-02 lute = -1.276501260e-07 pute = 2.775557562e-29
+ ua1 = 2.347446004e-09 lua1 = -5.120192258e-16
+ ub1 = -1.648087403e-18 lub1 = 4.244138946e-25
+ uc1 = -7.633649884e-11 luc1 = 4.487143608e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.196 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = 3.675e-10
+ vth0 = {-1.062772+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.85164386
+ k2 = -0.137927
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.66213569
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.35052697+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {3.1741044+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.49
+ etab = -6.25e-6
+ u0 = 0.0042057
+ ua = -2.005353e-9
+ ub = 2.0055289e-18
+ uc = 2.58041e-13
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 111898.0
+ a0 = 1.166315
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.45249595
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.028218739
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.82665932
+ pdiblc1 = 0.18776805
+ pdiblc2 = 0.0066944085
+ pdiblcb = -0.225
+ drout = 0.9981043
+ pscbe1 = 799968550.0
+ pscbe2 = 9.3174823e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.0852145
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.9262738e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.5675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.54112
+ kt2 = -0.042333
+ at = 105041.0
+ ute = -0.42503
+ ua1 = 2.9333e-10
+ ub1 = 5.4574e-20
+ uc1 = -5.8335e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.197 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.9635*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.3156e-8
+ lint = -8.1325e-9
+ vth0 = {9.612074778e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.972363322e-07 wvth0 = -8.993117806e-07 pvth0 = 1.765034266e-13
+ k1 = -1.820663869e+00 lk1 = 5.244804765e-07 wk1 = 8.949482650e-07 pk1 = -1.756470212e-13
+ k2 = 1.570841132e-03 lk2 = -2.737854379e-08 wk2 = 8.815870511e-08 pk2 = -1.730246826e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.812528741e+00 ldsub = -1.207106892e-06 wdsub = -2.311512125e-06 pdsub = 4.536689273e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {3.991766327e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.522401940e-07 wvoff = -1.888280002e-06 pvoff = 3.706032746e-13
+ nfactor = {-1.035637660e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.655559853e-06 wnfactor = 5.453341069e-06 pnfactor = -1.070299985e-12
+ eta0 = 8.304765258e+00 leta0 = -1.533764903e-06 weta0 = -3.487823512e-06 peta0 = 6.845376816e-13
+ etab = 4.529799288e-01 letab = -8.890533237e-08 wetab = -2.006426673e-07 petab = 3.937913310e-14
+ u0 = -4.022000678e-02 lu0 = 8.719211341e-09 wu0 = 1.897757190e-08 pu0 = -3.724633148e-15
+ ua = -3.838169482e-09 lua = 3.597177269e-16 wua = 7.018188546e-16 pua = -1.377424775e-22
+ ub = -6.681557303e-18 lub = 1.704970974e-24 wub = 3.768851024e-24 pub = -7.396935462e-31
+ uc = -3.838682792e-10 luc = 7.539055223e-17 wuc = 2.194742047e-16 puc = -4.307510479e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.212857852e+06 lvsat = -4.123448854e-01 wvsat = -8.483246505e-01 pvsat = 1.664964375e-7
+ a0 = 1.849664763e+00 la0 = -1.341176413e-07 wa0 = 9.408658508e-08 pa0 = -1.846590362e-14
+ ags = 1.249999985e+00 lags = 2.930155674e-15 wags = 6.663256613e-15 pags = -1.307763675e-21
+ a1 = 0.0
+ a2 = -8.824942107e+00 la2 = 1.820836380e-06 wa2 = 3.691368309e-06 pa2 = -7.244864011e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.583060888e+00 lketa = 3.051610943e-07 wketa = 6.667810102e-07 pketa = -1.308657750e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.014970397e+00 lpclm = -2.332238735e-07 wpclm = -3.048570274e-08 ppclm = 5.983276449e-15
+ pdiblc1 = 9.939370838e-02 lpdiblc1 = 1.734479016e-08 wpdiblc1 = 1.000998774e-07 ppdiblc1 = -1.964610244e-14
+ pdiblc2 = 6.397470244e-02 lpdiblc2 = -1.124211689e-08 wpdiblc2 = -1.817250159e-08 ppdiblc2 = 3.566626025e-15
+ pdiblcb = -9.722820553e+00 lpdiblcb = 1.864089751e-06 wpdiblcb = 4.934673143e-06 ppdiblcb = -9.685036244e-13
+ drout = 9.875979995e-01 ldrout = 2.062019073e-09 wdrout = 6.774321548e-15 pdrout = -1.329562238e-21
+ pscbe1 = 1.293148691e+09 lpscbe1 = -9.679400029e+01 wpscbe1 = -2.201889440e+02 ppscbe1 = 4.321538309e-5
+ pscbe2 = 1.583191728e-08 lpscbe2 = -1.278555580e-15 wpscbe2 = -3.288925542e-15 ppscbe2 = 6.455009714e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.297034939e+01 lbeta0 = -2.725166000e-06 wbeta0 = -4.457550399e-06 pbeta0 = 8.748611290e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.515150809e-07 lagidl = 3.031143249e-14 wagidl = 6.592771690e-14 pagidl = -1.293930336e-20
+ bgidl = 1.000000010e+09 lbgidl = -2.039252281e-06 wbgidl = -4.637317657e-06 pbgidl = 9.101424217e-13
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 1.0675e-9
+ dwc = -2.252e-8
+ xpart = 0.0
+ cgso = 5.47296e-11
+ cgdo = 5.47296e-11
+ cgbo = 0.0
+ cgdl = 6.932416e-12
+ cgsl = 6.932416e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.0006938237703
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 8.8756087e-11
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.37179002e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 6.379164807e-01 lkt1 = -2.314035949e-07 wkt1 = -5.731658334e-07 pkt1 = 1.124923923e-13
+ kt2 = 1.131417442e+00 lkt2 = -2.303661305e-07 wkt2 = -5.079194445e-07 pkt2 = 9.968680977e-14
+ at = 4.302022427e+03 lat = 1.977153543e-02 wat = 2.128918125e-01 pat = -4.178321157e-8
+ ute = -1.876135489e+00 lute = 2.848012187e-07 wute = -4.365889872e-15 pute = 8.568714627e-22
+ ua1 = -1.881882971e-10 lua1 = 9.450518858e-17 wua1 = -1.146674951e-15 pua1 = 2.250521593e-22
+ ub1 = 4.304954223e-18 lub1 = -8.342008745e-25 wub1 = -2.049391172e-25 pub1 = 4.022237583e-32
+ uc1 = -9.841078859e-10 luc1 = 1.816968155e-16 wuc1 = 4.736713851e-16 puc1 = -9.296511440e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
.ends sky130_fd_pr__pfet_01v8_hvt
* Well Proximity Effect Parameters
