* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 52
.param
+ sky130_fd_pr__pfet_01v8__toxe_mult = 1.0
+ sky130_fd_pr__pfet_01v8__rshp_mult = 1.0
+ sky130_fd_pr__pfet_01v8__overlap_mult = 9.5435e-1
+ sky130_fd_pr__pfet_01v8__ajunction_mult = 9.9626e-1
+ sky130_fd_pr__pfet_01v8__pjunction_mult = 1.0009e+0
+ sky130_fd_pr__pfet_01v8__lint_diff = 0.0
+ sky130_fd_pr__pfet_01v8__wint_diff = 0.0
+ sky130_fd_pr__pfet_01v8__dlc_diff = 0.0
+ sky130_fd_pr__pfet_01v8__dwc_diff = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 000, W = 1.26u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_0 = 0.66078
+ sky130_fd_pr__pfet_01v8__vsat_diff_0 = 16431.0
+ sky130_fd_pr__pfet_01v8__a0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_0 = -1.0309e-11
+ sky130_fd_pr__pfet_01v8__keta_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_0 = -0.019468
+ sky130_fd_pr__pfet_01v8__vth0_diff_0 = 0.035953
+ sky130_fd_pr__pfet_01v8__pditsd_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_0 = 0.00038997
+ sky130_fd_pr__pfet_01v8__b1_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_0 = -0.11598
+ sky130_fd_pr__pfet_01v8__ags_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_0 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_0 = 2.3766e-19
*
* sky130_fd_pr__pfet_01v8, Bin 001, W = 1.68u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_1 = 1.9928e-19
+ sky130_fd_pr__pfet_01v8__agidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_1 = 0.79871
+ sky130_fd_pr__pfet_01v8__vsat_diff_1 = -375.82
+ sky130_fd_pr__pfet_01v8__a0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_1 = -2.9528e-11
+ sky130_fd_pr__pfet_01v8__keta_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_1 = -0.023277
+ sky130_fd_pr__pfet_01v8__vth0_diff_1 = -0.017006
+ sky130_fd_pr__pfet_01v8__pditsd_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_1 = 0.00034579
+ sky130_fd_pr__pfet_01v8__b1_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_1 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_1 = -0.10952
+ sky130_fd_pr__pfet_01v8__ags_diff_1 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 002, W = 1.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_2 = -0.065739
+ sky130_fd_pr__pfet_01v8__ags_diff_2 = 0.081917
+ sky130_fd_pr__pfet_01v8__bgidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_2 = 3.0975e-19
+ sky130_fd_pr__pfet_01v8__agidl_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_2 = -0.079944
+ sky130_fd_pr__pfet_01v8__vsat_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_2 = -0.08023
+ sky130_fd_pr__pfet_01v8__pdits_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_2 = -1.8999e-11
+ sky130_fd_pr__pfet_01v8__keta_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_2 = -0.010076
+ sky130_fd_pr__pfet_01v8__vth0_diff_2 = -0.0058045
+ sky130_fd_pr__pfet_01v8__pditsd_diff_2 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_2 = 0.0014218
+ sky130_fd_pr__pfet_01v8__b1_diff_2 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 003, W = 1.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__b1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_3 = -0.068427
+ sky130_fd_pr__pfet_01v8__ags_diff_3 = 0.061544
+ sky130_fd_pr__pfet_01v8__bgidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_3 = 3.4961e-19
+ sky130_fd_pr__pfet_01v8__nfactor_diff_3 = 0.074091
+ sky130_fd_pr__pfet_01v8__vsat_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_3 = -0.070384
+ sky130_fd_pr__pfet_01v8__pdits_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_3 = -8.1128e-12
+ sky130_fd_pr__pfet_01v8__keta_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_3 = -0.013508
+ sky130_fd_pr__pfet_01v8__vth0_diff_3 = -0.00072299
+ sky130_fd_pr__pfet_01v8__pditsd_diff_3 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_3 = 0.0015782
*
* sky130_fd_pr__pfet_01v8, Bin 004, W = 1.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_4 = 0.0015543
+ sky130_fd_pr__pfet_01v8__vth0_diff_4 = -0.013035
+ sky130_fd_pr__pfet_01v8__b1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__cgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_4 = -0.066359
+ sky130_fd_pr__pfet_01v8__ags_diff_4 = 0.042979
+ sky130_fd_pr__pfet_01v8__ub_diff_4 = 3.2388e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_4 = 0.065236
+ sky130_fd_pr__pfet_01v8__vsat_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_4 = -0.044363
+ sky130_fd_pr__pfet_01v8__pdits_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_4 = -7.8248e-12
+ sky130_fd_pr__pfet_01v8__keta_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_4 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_4 = -0.014149
*
* sky130_fd_pr__pfet_01v8, Bin 005, W = 1.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__keta_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_5 = -0.01529
+ sky130_fd_pr__pfet_01v8__pditsd_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_5 = 0.0014113
+ sky130_fd_pr__pfet_01v8__vth0_diff_5 = -0.023687
+ sky130_fd_pr__pfet_01v8__b1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_5 = -0.073497
+ sky130_fd_pr__pfet_01v8__cgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_5 = 0.085625
+ sky130_fd_pr__pfet_01v8__ub_diff_5 = 3.2181e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_5 = 0.086719
+ sky130_fd_pr__pfet_01v8__vsat_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_5 = -0.081585
+ sky130_fd_pr__pfet_01v8__pdits_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_5 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_5 = -2.3572e-11
+ sky130_fd_pr__pfet_01v8__rdsw_diff_5 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 006, W = 1.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_6 = -0.025848
+ sky130_fd_pr__pfet_01v8__pditsd_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_6 = 0.00044436
+ sky130_fd_pr__pfet_01v8__vth0_diff_6 = -0.052157
+ sky130_fd_pr__pfet_01v8__b1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_6 = -0.10545
+ sky130_fd_pr__pfet_01v8__cgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_6 = 2.1528e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_6 = 0.84253
+ sky130_fd_pr__pfet_01v8__vsat_diff_6 = 110.49
+ sky130_fd_pr__pfet_01v8__agidl_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_6 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_6 = -2.6963e-11
*
* sky130_fd_pr__pfet_01v8, Bin 007, W = 1.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_7 = -2.9267e-11
+ sky130_fd_pr__pfet_01v8__rdsw_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_7 = -0.018493
+ sky130_fd_pr__pfet_01v8__pditsd_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_7 = 0.00020057
+ sky130_fd_pr__pfet_01v8__vth0_diff_7 = -0.036465
+ sky130_fd_pr__pfet_01v8__b1_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_7 = -0.12452
+ sky130_fd_pr__pfet_01v8__cgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_7 = 1.8997e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_7 = 0.41757
+ sky130_fd_pr__pfet_01v8__vsat_diff_7 = 20296.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_7 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_7 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 008, W = 1.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_8 = -2.1298e-11
+ sky130_fd_pr__pfet_01v8__rdsw_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_8 = -0.0092316
+ sky130_fd_pr__pfet_01v8__pditsd_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_8 = -0.00054138
+ sky130_fd_pr__pfet_01v8__vth0_diff_8 = 0.020532
+ sky130_fd_pr__pfet_01v8__b1_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_8 = -0.070563
+ sky130_fd_pr__pfet_01v8__cgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_8 = 1.5069e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_8 = -0.027492
+ sky130_fd_pr__pfet_01v8__vsat_diff_8 = 52497.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__pdits_diff_8 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_8 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 009, W = 1.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_9 = -7.015e-12
+ sky130_fd_pr__pfet_01v8__rdsw_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_9 = -0.01065
+ sky130_fd_pr__pfet_01v8__pditsd_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_9 = 0.00079381
+ sky130_fd_pr__pfet_01v8__vth0_diff_9 = 0.020733
+ sky130_fd_pr__pfet_01v8__b1_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_9 = -0.056914
+ sky130_fd_pr__pfet_01v8__cgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_9 = 2.4247e-19
+ sky130_fd_pr__pfet_01v8__bgidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_9 = -0.0015401
+ sky130_fd_pr__pfet_01v8__vsat_diff_9 = 15928.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_9 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_9 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 010, W = 2.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_10 = 4498.1
+ sky130_fd_pr__pfet_01v8__u0_diff_10 = 0.00042911
+ sky130_fd_pr__pfet_01v8__vth0_diff_10 = -0.052739
+ sky130_fd_pr__pfet_01v8__cgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_10 = -2.6742e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_10 = 0.88313
+ sky130_fd_pr__pfet_01v8__ub_diff_10 = 2.047e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_10 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_10 = -0.018259
+ sky130_fd_pr__pfet_01v8__voff_diff_10 = -0.13233
+ sky130_fd_pr__pfet_01v8__a0_diff_10 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 011, W = 3.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_11 = -0.055855
+ sky130_fd_pr__pfet_01v8__a0_diff_11 = -0.087355
+ sky130_fd_pr__pfet_01v8__pditsd_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_11 = 26714.0
+ sky130_fd_pr__pfet_01v8__u0_diff_11 = 0.0013928
+ sky130_fd_pr__pfet_01v8__vth0_diff_11 = -0.014131
+ sky130_fd_pr__pfet_01v8__cgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_11 = -3.8e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_11 = -0.025198
+ sky130_fd_pr__pfet_01v8__ub_diff_11 = 3.7335e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_11 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_11 = 0.06717
+ sky130_fd_pr__pfet_01v8__k2_diff_11 = -0.015275
*
* sky130_fd_pr__pfet_01v8, Bin 012, W = 3.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_12 = 0.060238
+ sky130_fd_pr__pfet_01v8__k2_diff_12 = -0.010456
+ sky130_fd_pr__pfet_01v8__voff_diff_12 = -0.051762
+ sky130_fd_pr__pfet_01v8__a0_diff_12 = -0.072023
+ sky130_fd_pr__pfet_01v8__pditsd_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_12 = 0.0018113
+ sky130_fd_pr__pfet_01v8__vth0_diff_12 = -0.010181
+ sky130_fd_pr__pfet_01v8__cgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_12 = -7.0667e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_12 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_12 = 0.011369
+ sky130_fd_pr__pfet_01v8__ub_diff_12 = 3.9754e-19
*
* sky130_fd_pr__pfet_01v8, Bin 013, W = 3.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_13 = 0.046528
+ sky130_fd_pr__pfet_01v8__ub_diff_13 = 3.83e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_13 = 0.034881
+ sky130_fd_pr__pfet_01v8__k2_diff_13 = -0.0085688
+ sky130_fd_pr__pfet_01v8__voff_diff_13 = -0.048343
+ sky130_fd_pr__pfet_01v8__a0_diff_13 = -0.041037
+ sky130_fd_pr__pfet_01v8__eta0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_13 = 0.0017986
+ sky130_fd_pr__pfet_01v8__vsat_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_13 = -0.00035839
+ sky130_fd_pr__pfet_01v8__cgidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_13 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_13 = -2.9121e-12
*
* sky130_fd_pr__pfet_01v8, Bin 014, W = 3.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_14 = -4.0591e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_14 = 0.038794
+ sky130_fd_pr__pfet_01v8__ub_diff_14 = 4.1037e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_14 = 0.015787
+ sky130_fd_pr__pfet_01v8__k2_diff_14 = -0.008116
+ sky130_fd_pr__pfet_01v8__voff_diff_14 = -0.038421
+ sky130_fd_pr__pfet_01v8__eta0_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_14 = -0.020215
+ sky130_fd_pr__pfet_01v8__pditsd_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_14 = 0.0019509
+ sky130_fd_pr__pfet_01v8__vsat_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_14 = 0.0024235
+ sky130_fd_pr__pfet_01v8__cgidl_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_14 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_14 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 015, W = 3.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_15 = 5.2325e-13
+ sky130_fd_pr__pfet_01v8__bgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_15 = 0.84448
+ sky130_fd_pr__pfet_01v8__ub_diff_15 = 1.6415e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_15 = -0.019065
+ sky130_fd_pr__pfet_01v8__pdits_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_15 = -0.097102
+ sky130_fd_pr__pfet_01v8__eta0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_15 = 0.00044761
+ sky130_fd_pr__pfet_01v8__vsat_diff_15 = -7259.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_15 = -0.027484
+ sky130_fd_pr__pfet_01v8__cgidl_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_15 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_15 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 016, W = 3.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_16 = 2.0071e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_16 = 0.33097
+ sky130_fd_pr__pfet_01v8__tvoff_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_16 = 1.9453e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_16 = -0.015561
+ sky130_fd_pr__pfet_01v8__pdits_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_16 = -0.12118
+ sky130_fd_pr__pfet_01v8__eta0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_16 = 0.00055244
+ sky130_fd_pr__pfet_01v8__vsat_diff_16 = 8567.5
+ sky130_fd_pr__pfet_01v8__vth0_diff_16 = -0.0057243
+ sky130_fd_pr__pfet_01v8__cgidl_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_16 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_16 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 017, W = 3.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_17 = -0.057073
+ sky130_fd_pr__pfet_01v8__ua_diff_17 = -5.0889e-11
+ sky130_fd_pr__pfet_01v8__tvoff_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_17 = 2.6612e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_17 = -0.0073251
+ sky130_fd_pr__pfet_01v8__pdits_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_17 = -0.089917
+ sky130_fd_pr__pfet_01v8__eta0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_17 = 0.00020589
+ sky130_fd_pr__pfet_01v8__vsat_diff_17 = 56793.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_17 = -0.017796
+ sky130_fd_pr__pfet_01v8__cgidl_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_17 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_17 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 018, W = 3.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_18 = 0.13485
+ sky130_fd_pr__pfet_01v8__ua_diff_18 = 9.2994e-13
+ sky130_fd_pr__pfet_01v8__tvoff_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_18 = 2.2388e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_18 = -0.015495
+ sky130_fd_pr__pfet_01v8__pdits_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_18 = -0.058923
+ sky130_fd_pr__pfet_01v8__eta0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_18 = 0.00093426
+ sky130_fd_pr__pfet_01v8__vsat_diff_18 = 15986.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_18 = 0.0018784
+ sky130_fd_pr__pfet_01v8__cgidl_diff_18 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_18 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 019, W = 5.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_19 = -0.039041
+ sky130_fd_pr__pfet_01v8__ua_diff_19 = -9.3266e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_19 = 0.040564
+ sky130_fd_pr__pfet_01v8__ub_diff_19 = 2.6349e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_19 = -0.009616
+ sky130_fd_pr__pfet_01v8__pdits_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_19 = -0.038421
+ sky130_fd_pr__pfet_01v8__eta0_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_19 = -0.045026
+ sky130_fd_pr__pfet_01v8__pditsd_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_19 = 0.0010965
+ sky130_fd_pr__pfet_01v8__vsat_diff_19 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_19 = 0.0069
*
* sky130_fd_pr__pfet_01v8, Bin 020, W = 5.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__u0_diff_20 = 0.0012594
+ sky130_fd_pr__pfet_01v8__vth0_diff_20 = 0.0013777
+ sky130_fd_pr__pfet_01v8__cgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_20 = -3.626e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_20 = 0.048112
+ sky130_fd_pr__pfet_01v8__ub_diff_20 = 2.7353e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_20 = 0.034261
+ sky130_fd_pr__pfet_01v8__k2_diff_20 = -0.011931
+ sky130_fd_pr__pfet_01v8__voff_diff_20 = -0.043221
+ sky130_fd_pr__pfet_01v8__a0_diff_20 = -0.039782
+ sky130_fd_pr__pfet_01v8__pditsd_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_20 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_20 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 021, W = 5.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_21 = 0.0016298
+ sky130_fd_pr__pfet_01v8__vth0_diff_21 = 0.0048083
+ sky130_fd_pr__pfet_01v8__cgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_21 = -2.4508e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_21 = 0.056607
+ sky130_fd_pr__pfet_01v8__ub_diff_21 = 3.1849e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_21 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_21 = 0.011009
+ sky130_fd_pr__pfet_01v8__k2_diff_21 = -0.011887
+ sky130_fd_pr__pfet_01v8__voff_diff_21 = -0.043022
+ sky130_fd_pr__pfet_01v8__a0_diff_21 = -0.012854
*
* sky130_fd_pr__pfet_01v8, Bin 022, W = 5.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_22 = -0.041062
+ sky130_fd_pr__pfet_01v8__a0_diff_22 = -0.011503
+ sky130_fd_pr__pfet_01v8__pditsd_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_22 = 0.0017941
+ sky130_fd_pr__pfet_01v8__vth0_diff_22 = 0.00086421
+ sky130_fd_pr__pfet_01v8__cgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_22 = -2.9796e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_22 = 0.060845
+ sky130_fd_pr__pfet_01v8__ub_diff_22 = 3.5456e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_22 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_22 = 0.0099482
+ sky130_fd_pr__pfet_01v8__k2_diff_22 = -0.012109
*
* sky130_fd_pr__pfet_01v8, Bin 023, W = 5.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_23 = -0.014758
+ sky130_fd_pr__pfet_01v8__voff_diff_23 = -0.12628
+ sky130_fd_pr__pfet_01v8__a0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_23 = -2987.4
+ sky130_fd_pr__pfet_01v8__u0_diff_23 = 0.00044006
+ sky130_fd_pr__pfet_01v8__vth0_diff_23 = -0.025813
+ sky130_fd_pr__pfet_01v8__cgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_23 = -1.5205e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_23 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_23 = 0.59286
+ sky130_fd_pr__pfet_01v8__ub_diff_23 = 1.6711e-19
*
* sky130_fd_pr__pfet_01v8, Bin 024, W = 5.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_24 = 0.28414
+ sky130_fd_pr__pfet_01v8__ub_diff_24 = 1.6768e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_24 = -0.011236
+ sky130_fd_pr__pfet_01v8__voff_diff_24 = -0.099324
+ sky130_fd_pr__pfet_01v8__a0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_24 = 0.00032449
+ sky130_fd_pr__pfet_01v8__vsat_diff_24 = 15165.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_24 = -0.016291
+ sky130_fd_pr__pfet_01v8__cgidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_24 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_24 = -8.5792e-12
*
* sky130_fd_pr__pfet_01v8, Bin 025, W = 5.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_25 = -5.3917e-13
+ sky130_fd_pr__pfet_01v8__bgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_25 = 0.11082
+ sky130_fd_pr__pfet_01v8__ub_diff_25 = 2.4381e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_25 = -0.0081573
+ sky130_fd_pr__pfet_01v8__voff_diff_25 = -0.067969
+ sky130_fd_pr__pfet_01v8__eta0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_25 = 0.00060876
+ sky130_fd_pr__pfet_01v8__vsat_diff_25 = 7602.9
+ sky130_fd_pr__pfet_01v8__vth0_diff_25 = -0.02575
+ sky130_fd_pr__pfet_01v8__cgidl_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_25 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_25 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 026, W = 5.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_26 = 5.7453e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_26 = 0.17526
+ sky130_fd_pr__pfet_01v8__ub_diff_26 = 2.8055e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_26 = -0.015244
+ sky130_fd_pr__pfet_01v8__pdits_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_26 = -0.041918
+ sky130_fd_pr__pfet_01v8__eta0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_26 = 0.0012472
+ sky130_fd_pr__pfet_01v8__vsat_diff_26 = 7612.8
+ sky130_fd_pr__pfet_01v8__vth0_diff_26 = -0.0033941
+ sky130_fd_pr__pfet_01v8__cgidl_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_26 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_26 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 027, W = 7.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_27 = -1.0829e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_27 = -0.077875
+ sky130_fd_pr__pfet_01v8__tvoff_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_27 = 0.090396
+ sky130_fd_pr__pfet_01v8__ub_diff_27 = 2.9028e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_27 = -0.01015
+ sky130_fd_pr__pfet_01v8__pdits_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_27 = -0.031586
+ sky130_fd_pr__pfet_01v8__eta0_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_27 = -0.13471
+ sky130_fd_pr__pfet_01v8__pditsd_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_27 = 0.0012178
+ sky130_fd_pr__pfet_01v8__vsat_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_27 = -0.0010962
+ sky130_fd_pr__pfet_01v8__cgidl_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_27 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_27 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 028, W = 7.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_28 = 0.0037674
+ sky130_fd_pr__pfet_01v8__ua_diff_28 = -7.2465e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_28 = 0.057344
+ sky130_fd_pr__pfet_01v8__ub_diff_28 = 2.958e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_28 = -0.012893
+ sky130_fd_pr__pfet_01v8__pdits_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_28 = -0.043436
+ sky130_fd_pr__pfet_01v8__eta0_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_28 = -0.066733
+ sky130_fd_pr__pfet_01v8__pditsd_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_28 = 0.0014119
+ sky130_fd_pr__pfet_01v8__vsat_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_28 = 0.0035411
+ sky130_fd_pr__pfet_01v8__cgidl_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_28 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_28 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 029, W = 7.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__bgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_29 = 0.06067
+ sky130_fd_pr__pfet_01v8__ua_diff_29 = -3.5733e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_29 = 0.015769
+ sky130_fd_pr__pfet_01v8__ub_diff_29 = 3.6594e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_29 = -0.012367
+ sky130_fd_pr__pfet_01v8__pdits_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_29 = -0.045297
+ sky130_fd_pr__pfet_01v8__eta0_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_29 = -0.019174
+ sky130_fd_pr__pfet_01v8__pditsd_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_29 = 0.0018877
+ sky130_fd_pr__pfet_01v8__vsat_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_29 = 0.00080521
+ sky130_fd_pr__pfet_01v8__cgidl_diff_29 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_29 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 030, W = 7.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_30 = -5.0977e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_30 = 0.093465
+ sky130_fd_pr__pfet_01v8__ub_diff_30 = 3.9461e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_30 = -0.014248
+ sky130_fd_pr__pfet_01v8__k2_diff_30 = -0.01321
+ sky130_fd_pr__pfet_01v8__voff_diff_30 = -0.050926
+ sky130_fd_pr__pfet_01v8__a0_diff_30 = 0.01682
+ sky130_fd_pr__pfet_01v8__pditsd_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_30 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_30 = 0.0020367
+ sky130_fd_pr__pfet_01v8__vth0_diff_30 = -0.00025351
*
* sky130_fd_pr__pfet_01v8, Bin 031, W = 7.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__u0_diff_31 = 0.00036257
+ sky130_fd_pr__pfet_01v8__vth0_diff_31 = -0.027514
+ sky130_fd_pr__pfet_01v8__cgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_31 = -3.5805e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_31 = 0.57096
+ sky130_fd_pr__pfet_01v8__ub_diff_31 = 1.4685e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_31 = -0.017121
+ sky130_fd_pr__pfet_01v8__voff_diff_31 = -0.12723
+ sky130_fd_pr__pfet_01v8__a0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_31 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_31 = -4716.5
*
* sky130_fd_pr__pfet_01v8, Bin 032, W = 7.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_32 = 8570.6
+ sky130_fd_pr__pfet_01v8__u0_diff_32 = 0.00050926
+ sky130_fd_pr__pfet_01v8__vth0_diff_32 = -0.014703
+ sky130_fd_pr__pfet_01v8__cgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_32 = 4.8344e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_32 = 0.21159
+ sky130_fd_pr__pfet_01v8__ub_diff_32 = 1.885e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_32 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_32 = -0.014444
+ sky130_fd_pr__pfet_01v8__voff_diff_32 = -0.047262
+ sky130_fd_pr__pfet_01v8__a0_diff_32 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 033, W = 7.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_33 = -0.041527
+ sky130_fd_pr__pfet_01v8__a0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_33 = 11761.0
+ sky130_fd_pr__pfet_01v8__u0_diff_33 = 0.00061072
+ sky130_fd_pr__pfet_01v8__vth0_diff_33 = -0.023852
+ sky130_fd_pr__pfet_01v8__cgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_33 = 8.1783e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_33 = 0.10437
+ sky130_fd_pr__pfet_01v8__ub_diff_33 = 2.2026e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_33 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_33 = -0.010822
*
* sky130_fd_pr__pfet_01v8, Bin 034, W = 7.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_34 = -0.016
+ sky130_fd_pr__pfet_01v8__voff_diff_34 = -0.057579
+ sky130_fd_pr__pfet_01v8__a0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_34 = 2998.3
+ sky130_fd_pr__pfet_01v8__u0_diff_34 = 0.0013699
+ sky130_fd_pr__pfet_01v8__vth0_diff_34 = -0.0020103
+ sky130_fd_pr__pfet_01v8__cgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_34 = 1.2152e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_34 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_34 = 0.27919
+ sky130_fd_pr__pfet_01v8__ub_diff_34 = 2.8017e-19
*
* sky130_fd_pr__pfet_01v8, Bin 035, W = 0.42u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_35 = 0.23441
+ sky130_fd_pr__pfet_01v8__ub_diff_35 = 3.3494e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_35 = -0.0066897
+ sky130_fd_pr__pfet_01v8__voff_diff_35 = -0.095705
+ sky130_fd_pr__pfet_01v8__a0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_35 = 0.0017171
+ sky130_fd_pr__pfet_01v8__vsat_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_35 = -0.031999
+ sky130_fd_pr__pfet_01v8__cgidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_35 = -3.9603e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_35 = 9.6587e-10
+ sky130_fd_pr__pfet_01v8__agidl_diff_35 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_35 = -8.8177e-12
*
* sky130_fd_pr__pfet_01v8, Bin 036, W = 0.42u, L = 20.0u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_36 = 1.8701e-9
+ sky130_fd_pr__pfet_01v8__ua_diff_36 = -4.9955e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_36 = 0.029222
+ sky130_fd_pr__pfet_01v8__ub_diff_36 = 7.6707e-21
+ sky130_fd_pr__pfet_01v8__pdits_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_36 = 0.006486
+ sky130_fd_pr__pfet_01v8__voff_diff_36 = -0.030456
+ sky130_fd_pr__pfet_01v8__eta0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_36 = 0.00012895
+ sky130_fd_pr__pfet_01v8__vsat_diff_36 = 20004.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_36 = 0.002147
+ sky130_fd_pr__pfet_01v8__cgidl_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_36 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_36 = -7.3618e-8
*
* sky130_fd_pr__pfet_01v8, Bin 037, W = 0.42u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_37 = -7.1448e-10
+ sky130_fd_pr__pfet_01v8__agidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_37 = 7.9686e-10
+ sky130_fd_pr__pfet_01v8__ua_diff_37 = -4.996e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_37 = 0.051268
+ sky130_fd_pr__pfet_01v8__ub_diff_37 = -7.0453e-20
+ sky130_fd_pr__pfet_01v8__tvoff_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_37 = 0.0031615
+ sky130_fd_pr__pfet_01v8__pdits_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_37 = -0.037179
+ sky130_fd_pr__pfet_01v8__eta0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_37 = -0.00037323
+ sky130_fd_pr__pfet_01v8__vsat_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_37 = 0.022099
+ sky130_fd_pr__pfet_01v8__cgidl_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_37 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_37 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 038, W = 0.42u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_38 = -1.9909e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_38 = 1.7302e-10
+ sky130_fd_pr__pfet_01v8__ua_diff_38 = -4.9282e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_38 = 0.04431
+ sky130_fd_pr__pfet_01v8__tvoff_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_38 = 1.428e-20
+ sky130_fd_pr__pfet_01v8__k2_diff_38 = -0.001698
+ sky130_fd_pr__pfet_01v8__pdits_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_38 = -0.036994
+ sky130_fd_pr__pfet_01v8__eta0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_38 = 0.00044339
+ sky130_fd_pr__pfet_01v8__vsat_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_38 = 0.00056812
+ sky130_fd_pr__pfet_01v8__cgidl_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_38 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_38 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 039, W = 0.42u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_39 = 3.6214e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_39 = 3.3703e-9
+ sky130_fd_pr__pfet_01v8__bgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_39 = 0.01066
+ sky130_fd_pr__pfet_01v8__ua_diff_39 = -7.1907e-12
+ sky130_fd_pr__pfet_01v8__tvoff_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_39 = 1.4267e-20
+ sky130_fd_pr__pfet_01v8__k2_diff_39 = 0.0016675
+ sky130_fd_pr__pfet_01v8__pdits_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_39 = -0.030352
+ sky130_fd_pr__pfet_01v8__eta0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_39 = 0.00029384
+ sky130_fd_pr__pfet_01v8__vsat_diff_39 = 20019.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_39 = 0.0048275
+ sky130_fd_pr__pfet_01v8__cgidl_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_39 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_39 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 040, W = 0.42u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_40 = -5.0608e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_40 = 2.6414e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_40 = -2.7512e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_40 = 1.1081
+ sky130_fd_pr__pfet_01v8__ub_diff_40 = 2.1195e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_40 = -0.030116
+ sky130_fd_pr__pfet_01v8__voff_diff_40 = -0.10278
+ sky130_fd_pr__pfet_01v8__a0_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_40 = 19687.0
+ sky130_fd_pr__pfet_01v8__u0_diff_40 = 0.00034139
+ sky130_fd_pr__pfet_01v8__vth0_diff_40 = 0.021587
+ sky130_fd_pr__pfet_01v8__cgidl_diff_40 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_40 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 041, W = 0.42u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__cgidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_41 = -7.5986e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_41 = 7.2273e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_41 = -2.732e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_41 = 1.1484
+ sky130_fd_pr__pfet_01v8__ub_diff_41 = 2.7027e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_41 = -0.023178
+ sky130_fd_pr__pfet_01v8__voff_diff_41 = -0.19428
+ sky130_fd_pr__pfet_01v8__a0_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_41 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_41 = 19660.0
+ sky130_fd_pr__pfet_01v8__u0_diff_41 = 0.00049786
+ sky130_fd_pr__pfet_01v8__vth0_diff_41 = 0.039021
*
* sky130_fd_pr__pfet_01v8, Bin 042, W = 0.42u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__u0_diff_42 = 0.0011703
+ sky130_fd_pr__pfet_01v8__vth0_diff_42 = -0.017565
+ sky130_fd_pr__pfet_01v8__cgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_42 = -4.3583e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_42 = 4.4592e-9
+ sky130_fd_pr__pfet_01v8__agidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_42 = -1.505e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_42 = 0.14181
+ sky130_fd_pr__pfet_01v8__ub_diff_42 = 2.7814e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_42 = -0.0065428
+ sky130_fd_pr__pfet_01v8__voff_diff_42 = -0.089
+ sky130_fd_pr__pfet_01v8__a0_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_42 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_42 = 20466.0
*
* sky130_fd_pr__pfet_01v8, Bin 043, W = 0.55u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pditsd_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_43 = 20224.0
+ sky130_fd_pr__pfet_01v8__u0_diff_43 = 0.0011785
+ sky130_fd_pr__pfet_01v8__vth0_diff_43 = -0.038893
+ sky130_fd_pr__pfet_01v8__cgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_43 = -3.9087e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_43 = -5.0176e-11
+ sky130_fd_pr__pfet_01v8__agidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_43 = -3.0087e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_43 = 0.14077
+ sky130_fd_pr__pfet_01v8__ub_diff_43 = 2.7797e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_43 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_43 = -0.01132
+ sky130_fd_pr__pfet_01v8__voff_diff_43 = -0.083804
+ sky130_fd_pr__pfet_01v8__a0_diff_43 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 044, W = 0.55u, L = 2.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__voff_diff_44 = -0.071307
+ sky130_fd_pr__pfet_01v8__a0_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_44 = 0.001722
+ sky130_fd_pr__pfet_01v8__vth0_diff_44 = 0.00059536
+ sky130_fd_pr__pfet_01v8__cgidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_44 = -7.4675e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_44 = 2.2895e-10
+ sky130_fd_pr__pfet_01v8__agidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_44 = -1.7426e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_44 = 0.10072
+ sky130_fd_pr__pfet_01v8__ub_diff_44 = 3.4467e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_44 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_44 = -0.0083627
*
* sky130_fd_pr__pfet_01v8, Bin 045, W = 0.55u, L = 4.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__pdits_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_45 = 0.00078773
+ sky130_fd_pr__pfet_01v8__voff_diff_45 = -0.035423
+ sky130_fd_pr__pfet_01v8__a0_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_45 = 20043.0
+ sky130_fd_pr__pfet_01v8__u0_diff_45 = 9.6015e-5
+ sky130_fd_pr__pfet_01v8__vth0_diff_45 = 0.0055575
+ sky130_fd_pr__pfet_01v8__cgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_45 = 1.6912e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_45 = 1.5334e-10
+ sky130_fd_pr__pfet_01v8__agidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_45 = -4.8743e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_45 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_45 = 0.029362
+ sky130_fd_pr__pfet_01v8__ub_diff_45 = -1.3062e-20
*
* sky130_fd_pr__pfet_01v8, Bin 046, W = 0.55u, L = 8.0u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__bgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_46 = 0.1837
+ sky130_fd_pr__pfet_01v8__ub_diff_46 = 3.1309e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_46 = -0.011371
+ sky130_fd_pr__pfet_01v8__voff_diff_46 = -0.082567
+ sky130_fd_pr__pfet_01v8__a0_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_46 = 0.0016571
+ sky130_fd_pr__pfet_01v8__vsat_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_46 = -0.021094
+ sky130_fd_pr__pfet_01v8__cgidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_46 = -7.5216e-8
+ sky130_fd_pr__pfet_01v8__b1_diff_46 = -1.295e-11
+ sky130_fd_pr__pfet_01v8__agidl_diff_46 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_46 = -7.5875e-12
*
* sky130_fd_pr__pfet_01v8, Bin 047, W = 0.55u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__agidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_47 = 2.5223e-9
+ sky130_fd_pr__pfet_01v8__ua_diff_47 = -2.3128e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_47 = 1.0026
+ sky130_fd_pr__pfet_01v8__ub_diff_47 = 2.367e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_47 = -0.024865
+ sky130_fd_pr__pfet_01v8__voff_diff_47 = -0.1571
+ sky130_fd_pr__pfet_01v8__eta0_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_47 = 0.00026524
+ sky130_fd_pr__pfet_01v8__vsat_diff_47 = 20030.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_47 = 0.029647
+ sky130_fd_pr__pfet_01v8__cgidl_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_47 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_47 = 2.6947e-8
*
* sky130_fd_pr__pfet_01v8, Bin 048, W = 0.55u, L = 0.5u
* ----------------------------------
+ sky130_fd_pr__pfet_01v8__b0_diff_48 = -6.8221e-8
+ sky130_fd_pr__pfet_01v8__agidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_48 = 3.3139e-10
+ sky130_fd_pr__pfet_01v8__ua_diff_48 = -1.2629e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_48 = 0.10376
+ sky130_fd_pr__pfet_01v8__ub_diff_48 = 2.9391e-19
+ sky130_fd_pr__pfet_01v8__tvoff_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_48 = -0.018886
+ sky130_fd_pr__pfet_01v8__pdits_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_48 = -0.080025
+ sky130_fd_pr__pfet_01v8__eta0_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_48 = 0.0011564
+ sky130_fd_pr__pfet_01v8__vsat_diff_48 = 20219.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_48 = -0.0020992
+ sky130_fd_pr__pfet_01v8__cgidl_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_48 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_48 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 049, W = 0.64u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__pclm_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_49 = 1.3673e-7
+ sky130_fd_pr__pfet_01v8__agidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_49 = 6.4955e-10
+ sky130_fd_pr__pfet_01v8__ua_diff_49 = -1.2078e-10
+ sky130_fd_pr__pfet_01v8__bgidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_49 = 1.0867
+ sky130_fd_pr__pfet_01v8__tvoff_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__ub_diff_49 = 2.2638e-19
+ sky130_fd_pr__pfet_01v8__k2_diff_49 = -0.013115
+ sky130_fd_pr__pfet_01v8__pdits_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__voff_diff_49 = -0.005274
+ sky130_fd_pr__pfet_01v8__eta0_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__a0_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__u0_diff_49 = 3.2751e-5
+ sky130_fd_pr__pfet_01v8__vsat_diff_49 = 21578.0
+ sky130_fd_pr__pfet_01v8__vth0_diff_49 = -0.045409
+ sky130_fd_pr__pfet_01v8__cgidl_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_49 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_49 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 050, W = 0.84u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__kt1_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_50 = -2.4518e-11
+ sky130_fd_pr__pfet_01v8__bgidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_50 = 0.94934
+ sky130_fd_pr__pfet_01v8__ub_diff_50 = 2.7121e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_50 = -0.040295
+ sky130_fd_pr__pfet_01v8__voff_diff_50 = -0.04981
+ sky130_fd_pr__pfet_01v8__a0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_50 = -26.109
+ sky130_fd_pr__pfet_01v8__u0_diff_50 = 0.00057771
+ sky130_fd_pr__pfet_01v8__vth0_diff_50 = -0.042662
+ sky130_fd_pr__pfet_01v8__cgidl_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_50 = 0.0
+ sky130_fd_pr__pfet_01v8__rdsw_diff_50 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 051, W = 1.65u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__pfet_01v8__rdsw_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__kt1_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__pclm_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__b0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__b1_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__agidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__ua_diff_51 = -6.7472e-12
+ sky130_fd_pr__pfet_01v8__bgidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__nfactor_diff_51 = 0.52474
+ sky130_fd_pr__pfet_01v8__ub_diff_51 = 2.3163e-19
+ sky130_fd_pr__pfet_01v8__pdits_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__tvoff_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__ags_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__k2_diff_51 = -0.030703
+ sky130_fd_pr__pfet_01v8__voff_diff_51 = -0.081386
+ sky130_fd_pr__pfet_01v8__a0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__pditsd_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__eta0_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__vsat_diff_51 = 2387.5
+ sky130_fd_pr__pfet_01v8__u0_diff_51 = 0.0005622
+ sky130_fd_pr__pfet_01v8__vth0_diff_51 = 0.0012633
+ sky130_fd_pr__pfet_01v8__cgidl_diff_51 = 0.0
+ sky130_fd_pr__pfet_01v8__keta_diff_51 = 0.0
*
* sky130_fd_pr__pfet_01v8, Bin 052, W = 0.42u, L = 0.17u
* sky130_fd_pr__pfet_01v8, Bin 053, W = 0.55u, L = 0.18u
* sky130_fd_pr__pfet_01v8, Bin 054, W = 0.55u, L = 0.17u
* sky130_fd_pr__pfet_01v8, Bin 055, W = 0.64u, L = 0.17u
* sky130_fd_pr__pfet_01v8, Bin 056, W = 0.64u, L = 0.18u
* sky130_fd_pr__pfet_01v8, Bin 057, W = 0.84u, L = 0.18u
* sky130_fd_pr__pfet_01v8, Bin 058, W = 0.84u, L = 0.17u
* sky130_fd_pr__pfet_01v8, Bin 059, W = 1.12u, L = 0.18u
* sky130_fd_pr__pfet_01v8, Bin 060, W = 1.26u, L = 0.18u
* sky130_fd_pr__pfet_01v8, Bin 061, W = 1.00u, L = 0.17u
* sky130_fd_pr__pfet_01v8, Bin 062, W = 1.12u, L = 0.17u
* sky130_fd_pr__pfet_01v8, Bin 063, W = 1.68u, L = 0.18u
* sky130_fd_pr__pfet_01v8, Bin 064, W = 2.00u, L = 0.18u
* sky130_fd_pr__pfet_01v8, Bin 065, W = 1.12u, L = 0.15u
* -----------------------------------
.include "sky130_fd_pr_models/cells/sky130_fd_pr__pfet_01v8.pm3.spice"
