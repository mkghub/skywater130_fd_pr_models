* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 38
.param
+ sky130_fd_pr__nfet_01v8_lvt__toxe_mult = 0.948
+ sky130_fd_pr__nfet_01v8_lvt__rshn_mult = 1.0
+ sky130_fd_pr__nfet_01v8_lvt__overlap_mult = 0.86067
+ sky130_fd_pr__nfet_01v8_lvt__ajunction_mult = 0.82447
+ sky130_fd_pr__nfet_01v8_lvt__pjunction_mult = 0.75
+ sky130_fd_pr__nfet_01v8_lvt__lint_diff = 1.7325e-8
+ sky130_fd_pr__nfet_01v8_lvt__wint_diff = -3.2175e-8
+ sky130_fd_pr__nfet_01v8_lvt__dlc_diff = 1.1336e-8
+ sky130_fd_pr__nfet_01v8_lvt__dwc_diff = -3.2175e-8
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 000, W = 1.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_0 = -0.11762
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_0 = 0.0081846
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_0 = 0.0011221
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_0 = -0.2
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_0 = 2.7218e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_0 = 3.8431e-19
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0 = 0.69693
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0 = -0.010063
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 001, W = 1.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_1 = -0.075108
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_1 = 0.0080507
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_1 = -0.16121
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_1 = -1.1838e-5
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_1 = 2.8356e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_1 = 2.6855e-19
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1 = 0.46688
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1 = -0.0097119
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 002, W = 1.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2 = -0.0049317
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_2 = 0.012804
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_2 = 0.010192
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_2 = -0.027026
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_2 = -0.00023333
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_2 = -4.0716e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_2 = 2.4704e-19
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2 = 0.74
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 003, W = 1.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3 = 1.5029
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3 = -0.085482
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_3 = 0.0504
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_3 = -0.0029143
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_3 = 2.99e-11
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3 = -40000.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_3 = 1.9717e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 004, W = 1.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4 = 1.5356
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4 = -0.10708
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_4 = 0.030667
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_4 = -0.0033249
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_4 = 1.4975e-11
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4 = -33009.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_4 = 9.1673e-20
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 005, W = 1.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_5 = 4.9257e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5 = 0.94557
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5 = -0.022141
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_5 = 0.012134
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_5 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_5 = 0.0013608
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_5 = 1.0925e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5 = -20000.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_5 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 006, W = 1.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_6 = 2.7039e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6 = 1.4368
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6 = -0.014763
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_6 = -0.0011301
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_6 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_6 = -0.00050123
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_6 = -1.4498e-12
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6 = -19315.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_6 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 007, W = 3.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_7 = 2.237e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7 = 0.77957
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7 = -0.00050334
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_7 = -0.062405
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_7 = 0.0033279
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_7 = -0.078248
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_7 = 0.00059112
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_7 = -3.0348e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 008, W = 3.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_8 = -0.061971
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_8 = -2.3628e-5
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_8 = 9.4746e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_8 = 1.7506e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8 = 0.37696
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8 = -0.0060049
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_8 = -0.040092
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_8 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_8 = 0.00064808
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 009, W = 3.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_9 = -0.023335
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_9 = -0.00038842
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_9 = -1.8365e-13
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_9 = 1.1976e-19
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9 = 0.41662
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9 = 0.0001567
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_9 = 0.0088493
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_9 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_9 = 0.0056151
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 010, W = 3.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_10 = 9.1989e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_10 = -1.5913e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_10 = -0.0038906
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10 = -32682.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10 = -0.11138
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10 = 1.4545
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_10 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_10 = 0.054715
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 011, W = 3.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_11 = 0.036624
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_11 = 4.043e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_11 = 1.7433e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_11 = -0.0014474
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11 = -22283.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11 = -0.082765
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11 = 1.1674
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 012, W = 3.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_12 = 0.017873
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_12 = -7.4481e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_12 = 4.9896e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_12 = 0.00021131
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12 = -15131.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12 = -0.029909
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12 = 0.9639
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_12 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_12 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 013, W = 3.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_13 = 0.012552
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_13 = 1.7628e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_13 = 2.2271e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_13 = -0.00084741
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13 = -12681.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13 = -0.010116
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13 = 1.2538
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_13 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_13 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 014, W = 5.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14 = 0.62815
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_14 = 0.002812
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_14 = 9.5412e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_14 = 1.9897e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_14 = -0.065447
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_14 = -0.09371
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_14 = 0.00022119
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14 = -0.0093128
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 015, W = 5.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15 = 0.0010127
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15 = 0.48677
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_15 = -0.0061278
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_15 = -5.7198e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_15 = 2.1734e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_15 = 0.0010625
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_15 = -0.0092625
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_15 = 0.00026915
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 016, W = 5.0u, L = 4.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_16 = -0.035853
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_16 = -0.00010032
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16 = -0.011405
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16 = 0.10165
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_16 = 0.0081435
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_16 = 1.1846e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_16 = 1.4143e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_16 = 0.004933
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 017, W = 5.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_17 = -0.0019594
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17 = -26495.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17 = -0.09687
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17 = 1.35
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_17 = 0.059013
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_17 = 5.5844e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_17 = 1.0731e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 018, W = 5.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_18 = -0.0022255
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18 = -25421.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18 = -0.065606
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18 = 1.2946
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_18 = 0.037119
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_18 = 4.7069e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_18 = 6.8941e-20
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 019, W = 5.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_19 = 3.6894e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_19 = -0.00074934
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19 = -19755.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19 = -0.036018
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19 = 0.73262
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_19 = 0.014685
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_19 = -2.4883e-11
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 020, W = 5.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_20 = -3.9165e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_20 = 2.3083e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_20 = -0.00023099
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20 = -9270.2
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20 = -0.012834
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20 = 1.2218
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_20 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_20 = 0.0015349
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 021, W = 7.0u, L = 1.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_21 = -2.5325e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_21 = 2.2719e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_21 = 0.018948
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_21 = 0.016513
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_21 = 0.0006107
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21 = -4.4035e-5
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21 = 0.76771
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_21 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_21 = -0.0052929
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 022, W = 7.0u, L = 2.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_22 = 0.007281
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_22 = 4.94e-15
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_22 = 1.709e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_22 = -0.0096289
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_22 = -0.029399
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_22 = 5.1709e-5
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22 = -0.005971
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22 = 0.45812
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 023, W = 7.0u, L = 8.0u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_23 = 0.0064536
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_23 = -1.5075e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_23 = 1.907e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_23 = 0.0008694
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_23 = 0.01967
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_23 = 0.00045513
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23 = -0.0046908
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23 = 0.31335
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_23 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_23 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 024, W = 7.0u, L = 0.15u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_24 = 0.058237
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_24 = 5.0139e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_24 = -1.347e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_24 = -0.0060241
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24 = -27273.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24 = -0.11108
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24 = 1.3376
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_24 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_24 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 025, W = 7.0u, L = 0.18u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25 = 1.2595
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_25 = 0.032673
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_25 = 1.2484e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_25 = -2.7509e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_25 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_25 = -0.0035292
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25 = -24107.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25 = -0.059801
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 026, W = 7.0u, L = 0.25u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26 = -0.024267
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26 = 0.69726
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_26 = 0.015591
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_26 = 2.3711e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_26 = 3.4661e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_26 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_26 = 0.00018708
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26 = -17553.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 027, W = 7.0u, L = 0.5u
* ---------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_27 = -0.00025306
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27 = -5519.2
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27 = -0.0062576
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27 = 0.97342
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_27 = 0.0037121
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_27 = -1.3023e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_27 = 1.9461e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_27 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 028, W = 0.42u, L = 1.0u
* ----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_28 = 0.0012314
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28 = -0.025962
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28 = 0.015295
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_28 = 1.9154e-7
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_28 = 1.9078e-9
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_28 = 0.0065995
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_28 = 2.1038e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_28 = 5.2387e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 029, W = 0.42u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_29 = -0.0032316
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29 = -43064.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29 = -0.16083
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29 = 1.6738
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_29 = 0.04922
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_29 = 4.2051e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_29 = 2.7257e-19
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 030, W = 0.42u, L = 0.18u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_30 = 7.8237e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_30 = -0.0026177
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30 = -38284.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30 = -0.13533
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30 = 1.6291
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_30 = 0.021285
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_30 = 3.7522e-11
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 031, W = 0.55u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_31 = 9.4623e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_31 = -3.1689e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_31 = -0.0037292
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31 = -50482.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31 = -0.18325
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31 = 2.3213
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_31 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_31 = 0.032738
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 032, W = 0.64u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_32 = 2.3172e-10
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_32 = -4.2095e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_32 = -0.0014643
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32 = -36597.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32 = -0.18077
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32 = 2.2437
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_32 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_32 = 0.033141
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 033, W = 0.84u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_33 = 0.032169
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_33 = 8.1829e-11
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_33 = -2.9805e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_33 = -0.0026455
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33 = -30414.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33 = -0.17173
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33 = 1.9708
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 034, W = 1.65u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_34 = 0.05002
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_34 = 8.6394e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_34 = -6.9165e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_34 = -0.0045403
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34 = -31996.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34 = -0.11639
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34 = 1.8011
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_34 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_34 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 035, W = 3.01u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_35 = 0.052812
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_35 = 1.0147e-12
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_35 = -5.2128e-20
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_35 = -0.0041733
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35 = -34265.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35 = -0.10525
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35 = 1.268
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_35 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_35 = 0.0
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 036, W = 5.05u, L = 0.15u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36 = 1.4418
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_36 = 0.059239
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_36 = 5.1438e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_36 = 1.8875e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_36 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_36 = -0.0023005
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36 = -26664.0
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36 = -0.094492
*
* sky130_fd_pr__nfet_01v8_lvt, Bin 037, W = 5.05u, L = 0.25u
* -----------------------------------
+ sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37 = -0.031305
+ sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37 = 0.86841
+ sky130_fd_pr__nfet_01v8_lvt__voff_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__b1_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__keta_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__k2_diff_37 = 0.01431
+ sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ua_diff_37 = 1.7269e-13
+ sky130_fd_pr__nfet_01v8_lvt__ub_diff_37 = 3.3705e-19
+ sky130_fd_pr__nfet_01v8_lvt__a0_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__ags_diff_37 = 0.0
+ sky130_fd_pr__nfet_01v8_lvt__u0_diff_37 = -0.00060631
+ sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37 = -18688.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_01v8_lvt.pm3.spice"
