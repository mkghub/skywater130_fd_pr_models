* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
* Number of bins: 11
.param
+ sky130_fd_pr__nfet_05v0_nvt__toxe_mult = 1.0365
+ sky130_fd_pr__nfet_05v0_nvt__rshn_mult = 1.0
+ sky130_fd_pr__nfet_05v0_nvt__overlap_mult = 1.1614
+ sky130_fd_pr__nfet_05v0_nvt__ajunction_mult = 1.2643e+0
+ sky130_fd_pr__nfet_05v0_nvt__pjunction_mult = 1.1856e+0
+ sky130_fd_pr__nfet_05v0_nvt__lint_diff = -1.21275e-8
+ sky130_fd_pr__nfet_05v0_nvt__wint_diff = 2.252e-8
+ sky130_fd_pr__nfet_05v0_nvt__dlc_diff = -3.0000e-8
+ sky130_fd_pr__nfet_05v0_nvt__dwc_diff = 2.252e-8
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 000, W = 10.0u, L = 2.0u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_0 = -0.032984
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_0 = 0.057763
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_0 = 7.2807e-5
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_0 = -0.0067973
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_0 = -2.376e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_0 = 0.021482
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_0 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_0 = 0.0047929
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_0 = -1.1063e-18
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 001, W = 10.0u, L = 4.0u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_1 = -1.119e-18
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_1 = 0.077833
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_1 = 0.027909
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_1 = -0.002922
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_1 = -0.0064693
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_1 = -2.2842e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_1 = 0.013709
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_1 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_1 = 0.0032394
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 002, W = 10.0u, L = 0.9u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_2 = -1.0808e-18
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_2 = -0.14696
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_2 = 0.0022692
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_2 = -0.0072977
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_2 = -2.3876e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_2 = 864.93
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_2 = 0.027939
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_2 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_2 = 0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 003, W = 1.0u, L = 25.0u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_3 = -1.1915e-11
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_3 = 0.0166
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_3 = -8.2319e-19
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_3 = 0.11551
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_3 = 0.00089555
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_3 = -0.0041127
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_3 = -0.0071709
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_3 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_3 = -0.0033311
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 004, W = 1.0u, L = 2.0u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_4 = -0.0078839
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_4 = 0.0084729
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_4 = -2.0087e-11
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_4 = 0.014055
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_4 = -1.1143e-18
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_4 = 0.10719
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_4 = 0.06314
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_4 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_4 = -0.0012356
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 005, W = 1.0u, L = 4.0u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_5 = 0.00058708
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_5 = -0.0088249
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_5 = 0.0067298
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_5 = -1.6502e-11
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_5 = 0.019503
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_5 = -1.075e-18
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_5 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_5 = 0.11267
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_5 = 0.088664
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_5 = 0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 006, W = 1.0u, L = 8.0u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_6 = 0.044119
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_6 = -0.0019442
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_6 = -0.0072188
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_6 = 0.00092262
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_6 = -1.3916e-11
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_6 = 0.0087222
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_6 = -9.064e-19
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_6 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_6 = 0.13457
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 007, W = 1.0u, L = 0.9u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_7 = -0.032084
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_7 = 0.00069292
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_7 = -0.0092302
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_7 = 0.0096456
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_7 = -1.9874e-11
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_7 = 288.71
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_7 = -1.0787e-18
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_7 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_7 = 0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 008, W = 0.42u, L = 1.0u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_8 = 0.041165
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_8 = 4.35e-8
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_8 = 0.00055638
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_8 = -0.010837
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_8 = -0.010299
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_8 = -2.8046e-12
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_8 = 3.3176e-10
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_8 = -7.4006e-19
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_8 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_8 = 0.0
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 009, W = 0.42u, L = 0.9u
* -------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_9 = 0.13133
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_9 = 0.0023042
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_9 = -0.01127
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_9 = 0.020187
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_9 = 4.2431e-12
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_9 = -4479.0
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_9 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_9 = -3.7969e-19
*
* sky130_fd_pr__nfet_05v0_nvt, Bin 010, W = 0.7u, L = 0.9u
* ------------------------------------
+ sky130_fd_pr__nfet_05v0_nvt__vsat_diff_10 = -1768.2
+ sky130_fd_pr__nfet_05v0_nvt__vth0_diff_10 = 0.013913
+ sky130_fd_pr__nfet_05v0_nvt__b0_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__keta_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__b1_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__kt1_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__pclm_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_10 = 0.0061791
+ sky130_fd_pr__nfet_05v0_nvt__ags_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__u0_diff_10 = -0.010406
+ sky130_fd_pr__nfet_05v0_nvt__pdits_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__k2_diff_10 = 0.00086128
+ sky130_fd_pr__nfet_05v0_nvt__ua_diff_10 = -1.3004e-11
+ sky130_fd_pr__nfet_05v0_nvt__eta0_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__ub_diff_10 = -8.7248e-19
+ sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__voff_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__a0_diff_10 = 0.0
+ sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_10 = 0.0
.include "sky130_fd_pr_models/cells/sky130_fd_pr__nfet_05v0_nvt.pm3.spice"
