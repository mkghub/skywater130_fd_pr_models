* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_01v8__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__voff_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__nfet_01v8 d g s b
+ 
.param  l = 1u w = 1u ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 nf = 1.0
msky130_fd_pr__nfet_01v8 d g s b sky130_fd_pr__nfet_01v8__model l = {l} w = {w} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} nf = {nf}
.model sky130_fd_pr__nfet_01v8__model.0 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.5160869+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.54086565
+ k2 = -0.026708291
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.68453
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0314621
+ ua = -7.5795907e-10
+ ub = 1.57049e-18
+ uc = 4.9242e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.369451
+ ags = 0.380025
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 2.1073424e-24
+ keta = -0.0087946
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.026316
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030734587
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 754674160.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31303
+ kt2 = -0.045313337
+ at = 140000.0
+ ute = -1.8134
+ ua1 = 3.7602e-10
+ ub1 = -6.3962e-19
+ uc1 = 1.5829713e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.1 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.5160869+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.54086565
+ k2 = -0.026708291
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.68453
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0314621
+ ua = -7.5795907e-10
+ ub = 1.57049e-18
+ uc = 4.9242e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.369451
+ ags = 0.380025
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 2.1073424e-24
+ keta = -0.0087946
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.026316
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030734587
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 754674160.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31303
+ kt2 = -0.045313337
+ at = 140000.0
+ ute = -1.8134
+ ua1 = 3.7602e-10
+ ub1 = -6.3962e-19
+ uc1 = 1.5829713e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.2 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.166909460e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.838883101e-09 wvth0 = -6.033932022e-08 pvth0 = 4.833653817e-13
+ k1 = 5.415453773e-01 lk1 = -5.445149777e-09 wk1 = -6.789927122e-08 pk1 = 5.439265313e-13
+ k2 = -2.711805592e-02 lk2 = 3.282539101e-09 wk2 = 4.093220973e-08 pk2 = -3.278991727e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.049996442e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.154547359e-09 wvoff = -2.686651451e-08 pvoff = 2.152218983e-13
+ nfactor = 2.686034709e+00 lnfactor = -1.205390299e-08 wnfactor = -1.503083041e-07 pnfactor = 1.204087658e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.142325993e-02 lu0 = 3.111395108e-10 wu0 = 3.879809903e-09 pu0 = -3.108032685e-14
+ ua = -7.575504764e-10 lua = -3.273155509e-18 wua = -4.081519935e-17 pua = 3.269618276e-22
+ ub = 1.564807772e-18 lub = 4.551910922e-26 wub = 5.676086919e-25 pub = -4.546991763e-30
+ uc = 4.877037585e-11 luc = 3.778080112e-18 wuc = 4.711144720e-17 puc = -3.773997217e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.361739852e+00 la0 = 6.177235391e-08 wa0 = 7.702814400e-07 pa0 = -6.170559776e-12
+ ags = 3.816712633e-01 lags = -1.318786275e-08 wags = -1.644484186e-07 pags = 1.317361089e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 1.950752899e-24 lb1 = 1.254404981e-30 wb1 = 1.564202776e-29 pb1 = -1.253049370e-34
+ keta = -8.288371258e-03 lketa = -4.055290119e-09 wketa = -5.056816706e-08 pketa = 4.050907648e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.798002168e-02 lpclm = -3.337615616e-07 wpclm = -4.161899621e-06 ppclm = 3.334008721e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.074731372e-03 lpdiblc2 = -1.019510186e-11 wpdiblc2 = -1.271296502e-10 ppdiblc2 = 1.018408422e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.580421702e+08 lpscbe1 = -2.698040880e+01 wpscbe1 = -3.364370440e+02 ppscbe1 = 2.695125162e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.131867870e-01 lkt1 = 1.255986929e-09 wkt1 = 1.566175415e-08 pkt1 = -1.254629609e-13
+ kt2 = -4.539666594e-02 lkt2 = 6.675302662e-10 wkt2 = 8.323888313e-09 pkt2 = -6.668088796e-14
+ at = 140000.0
+ ute = -1.816357404e+00 lute = 2.369112785e-08 wute = 2.954207655e-07 pute = -2.366552532e-12
+ ua1 = 3.613845672e-10 lua1 = 1.172413201e-16 wua1 = 1.461961658e-15 pua1 = -1.171146198e-20
+ ub1 = -6.204600368e-19 lub1 = -1.534863647e-25 wub1 = -1.913925738e-24 pub1 = 1.533204951e-29
+ uc1 = 1.690921780e-11 luc1 = -8.647681916e-18 wuc1 = -1.078338198e-16 puc1 = 8.638336539e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.3 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.071728966e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.333597610e-08 wvth0 = 7.402623097e-08 pvth0 = -5.554608993e-14
+ k1 = 5.302997219e-01 lk1 = 3.965876745e-08 wk1 = 1.367515665e-07 pk1 = -2.768841837e-13
+ k2 = -2.048316993e-02 lk2 = -2.332856876e-08 wk2 = -6.801314992e-08 pk2 = 1.090573506e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 5.376480639e-01 ldsub = 8.964883236e-08 wdsub = 2.232778080e-06 pdsub = -8.955195066e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.094655827e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.575737635e-08 wvoff = 5.573196081e-08 pvoff = -1.160629101e-13
+ nfactor = 2.666085505e+00 lnfactor = 6.795808584e-08 wnfactor = -1.912644030e-07 pnfactor = 1.368353806e-12
+ eta0 = 7.407673693e-02 leta0 = 2.375694058e-08 weta0 = 5.916861913e-07 peta0 = -2.373126692e-12
+ etab = -6.482185296e-02 letab = -2.076843965e-08 wetab = -5.172551119e-07 petab = 2.074599561e-12
+ u0 = 3.194993327e-02 lu0 = -1.801234574e-09 wu0 = 3.764492127e-09 pu0 = -3.061781193e-14
+ ua = -7.771556207e-10 lua = 7.535888247e-17 wua = 1.365337502e-15 pua = -5.312815741e-21
+ ub = 1.668742330e-18 lub = -3.713401575e-25 wub = -2.134683279e-24 pub = 6.291323040e-30
+ uc = 5.890739593e-11 luc = -3.687933810e-17 wuc = -3.280617428e-16 puc = 1.127339656e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.490798641e+00 la0 = -4.558548281e-07 wa0 = -1.699489791e-06 pa0 = 3.735164101e-12
+ ags = 3.647656614e-01 lags = 5.461688862e-08 wags = -7.007562172e-07 pags = 3.468376900e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 4.539228699e-24 lb1 = -9.127417519e-30 wb1 = -3.128405553e-29 pb1 = 6.290554088e-35
+ keta = -1.651832020e-02 lketa = 2.895327386e-08 wketa = 8.733344889e-08 pketa = -1.480031059e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.228164149e-01 lpclm = 2.436875115e-06 wpclm = 8.531224325e-06 ppclm = -1.756931660e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.181986903e-03 lpdiblc2 = -4.403740832e-10 wpdiblc2 = -1.256119770e-08 ppdiblc2 = 5.088879447e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.023678574e+08 lpscbe1 = 1.963173455e+02 wpscbe1 = 6.728740879e+02 ppscbe1 = -1.353005796e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.112536839e-01 lkt1 = -6.497275977e-09 wkt1 = 3.446901913e-08 pkt1 = -2.008948760e-13
+ kt2 = -4.402024159e-02 lkt2 = -4.853013239e-09 wkt2 = -1.654486044e-08 pkt2 = 3.306234138e-14
+ at = 1.381328683e+05 lat = 7.488665797e-03 wat = 1.865113957e-01 pat = -7.480572945e-7
+ ute = -1.757166309e+00 lute = -2.137116870e-07 wute = -1.620152226e-06 pute = 5.316400804e-12
+ ua1 = 6.261329075e-10 lua1 = -9.446076166e-16 wua1 = -5.203440883e-15 pua1 = 1.502204122e-20
+ ub1 = -9.508554259e-19 lub1 = 1.171658836e-24 wub1 = 5.193865106e-24 pub1 = -1.317577850e-29
+ uc1 = -4.824542424e-13 luc1 = 6.110659282e-17 wuc1 = 1.704269561e-16 puc1 = -2.522107706e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.4 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.256581141e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.833840380e-09 wvth0 = -1.440555601e-07 pvth0 = 3.829697225e-13
+ k1 = 5.525508708e-01 lk1 = -5.083531333e-09 wk1 = -2.534878473e-07 pk1 = 5.078037662e-13
+ k2 = -3.311163166e-02 lk2 = 2.064565301e-09 wk2 = 8.878661258e-08 pk2 = -2.062334167e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 5.822320387e-01 wdsub = -2.220801299e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.030312872e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.819384981e-09 wvoff = 1.380733451e-07 pvoff = -2.816338128e-13
+ nfactor = 2.691123862e+00 lnfactor = 1.761130745e-08 wnfactor = 1.364137978e-06 pnfactor = -1.759227527e-12
+ eta0 = 8.604364330e-02 leta0 = -3.059472010e-10 weta0 = -6.037112053e-07 peta0 = 3.056165700e-14
+ etab = -7.513627443e-02 letab = -2.834536917e-11 wetab = 5.130723758e-07 petab = 2.831473690e-15
+ u0 = 3.078800555e-02 lu0 = 5.351534303e-10 wu0 = 1.512308431e-08 pu0 = -5.345751007e-14
+ ua = -7.785201420e-10 lua = 7.810264280e-17 wua = 2.603165964e-15 pua = -7.801823884e-21
+ ub = 1.523558700e-18 lub = -7.940694862e-26 wub = -2.950677856e-24 pub = 7.932113512e-30
+ uc = 3.955982554e-11 luc = 2.024485577e-18 wuc = 3.331570204e-16 puc = -2.022297756e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.152059407e+04 lvsat = -3.057589258e-03 wvsat = -1.518950790e-01 pvsat = 3.054284983e-7
+ a0 = 1.249877415e+00 la0 = 2.858620026e-08 wa0 = 1.578181166e-06 pa0 = -2.855530773e-12
+ ags = 4.177671586e-01 lags = -5.195777995e-08 wags = -1.557031386e-06 pags = 5.190163022e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.984076421e-03 lketa = 9.781949960e-09 wketa = 4.996770669e-07 pketa = -9.771378803e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.765408299e-01 lpclm = 2.522435828e-08 wpclm = 1.046784548e-06 ppclm = -2.519709882e-12
+ pdiblc1 = 4.137574096e-01 lpdiblc1 = -4.777106666e-08 wpdiblc1 = -2.373173546e-06 ppdiblc1 = 4.771944142e-12
+ pdiblc2 = 2.902975442e-03 lpdiblc2 = 1.206582560e-10 wpdiblc2 = 1.874078111e-08 ppdiblc2 = -1.205278630e-14
+ pdiblcb = -2.314169863e-02 lpdiblcb = -3.736646369e-09 wpdiblcb = -1.856293136e-07 ppdiblcb = 3.732608250e-13
+ drout = 5.375281665e-01 ldrout = 4.518604815e-08 wdrout = 2.244754862e-06 pdrout = -4.513721650e-12
+ pscbe1 = 7.596311908e+08 lpscbe1 = 8.117303628e+01 wpscbe1 = 4.032518339e+03 ppscbe1 = -8.108531420e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.255049513e-07 lalpha0 = -3.931186189e-13 walpha0 = -1.952936730e-11 palpha0 = 3.926937835e-17
+ alpha1 = 8.525468078e-01 lalpha1 = -5.121085457e-09 walpha1 = -2.544055510e-07 palpha1 = 5.115551203e-13
+ beta0 = 1.406763974e+01 lbeta0 = -4.175190849e-07 wbeta0 = -2.074153492e-05 pbeta0 = 4.170678804e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.106429615e-01 lkt1 = -7.725308033e-09 wkt1 = -4.492178678e-07 pkt1 = 7.716959447e-13
+ kt2 = -4.493098135e-02 lkt2 = -3.021710482e-09 wkt2 = -1.502150554e-07 pkt2 = 3.018444980e-13
+ at = 1.379939085e+05 lat = 7.768084158e-03 wat = 2.003923556e-01 pat = -7.759689345e-7
+ ute = -1.801420659e+00 lute = -1.247256600e-07 wute = -5.172338457e-06 pute = 1.245908715e-11
+ ua1 = 2.851161315e-10 lua1 = -2.588958578e-16 wua1 = -1.059415188e-14 pua1 = 2.586160742e-20
+ ub1 = -4.357671071e-19 lub1 = 1.359264559e-25 wub1 = 5.393875348e-24 pub1 = -1.357795629e-29
+ uc1 = 3.136246856e-11 luc1 = -2.926732120e-18 wuc1 = -1.003963420e-16 puc1 = 2.923569259e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.5 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.171853786e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.730281984e-09 wvth0 = 6.264239100e-08 pvth0 = 1.740423273e-13
+ k1 = 5.402511595e-01 lk1 = 7.348844679e-09 wk1 = 9.882211729e-07 pk1 = -7.472983274e-13
+ k2 = -2.611597326e-02 lk2 = -5.006548271e-09 wk2 = -4.201058587e-07 pk2 = 3.081479688e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 9.216734667e-01 ldsub = -3.431026432e-07 wdsub = -5.514221115e-06 pdsub = 3.328942642e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.009799929e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.459654747e-10 wvoff = -3.942667057e-08 pvoff = -1.022192820e-13
+ nfactor = 2.651060692e+00 lnfactor = 5.810659875e-08 wnfactor = -1.378147636e-06 pnfactor = 1.012636380e-12
+ eta0 = 2.098785464e-01 leta0 = -1.254765336e-07 weta0 = -4.861098268e-06 peta0 = 4.333868896e-12
+ etab = -1.514243402e-01 letab = 7.708256352e-08 wetab = 1.041452527e-06 petab = -5.312477862e-13
+ u0 = 3.290551512e-02 lu0 = -1.605195596e-09 wu0 = -3.838977123e-08 pu0 = 6.325351285e-16
+ ua = -5.246086823e-10 lua = -1.785475059e-16 wua = -5.159390749e-15 pua = 4.445976670e-23
+ ub = 1.302653397e-18 lub = 1.438810395e-25 wub = 5.412114832e-24 pub = -5.208802570e-31
+ uc = 8.743480464e-12 luc = 3.317321575e-17 wuc = 2.052528342e-16 puc = -7.294601488e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.011565249e+04 lvsat = -1.637493983e-03 wvsat = -1.155275070e-02 pvsat = 1.635724376e-7
+ a0 = 1.285218759e+00 la0 = -7.136336130e-09 wa0 = -4.131210800e-06 pa0 = 2.915442695e-12
+ ags = 2.421556360e-01 lags = 1.255478885e-07 wags = 1.867376187e-06 pags = 1.728819788e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.552025509e-03 lketa = -8.677943660e-10 wketa = -7.420484664e-07 pketa = 2.779809047e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.430483739e-01 lpclm = -4.200053613e-08 wpclm = -2.752738181e-06 ppclm = 1.320794500e-12
+ pdiblc1 = 3.886654915e-01 lpdiblc1 = -2.240850714e-08 wpdiblc1 = 1.333066290e-07 ppdiblc1 = 2.238429072e-12
+ pdiblc2 = 1.088563979e-03 lpdiblc2 = 1.954639961e-09 wpdiblc2 = 2.427070621e-08 ppdiblc2 = -1.764235717e-14
+ pdiblcb = -2.871660273e-02 lpdiblcb = 1.898388643e-09 wpdiblcb = 3.712586273e-07 ppdiblcb = -1.896337092e-13
+ drout = 6.003068905e-01 ldrout = -1.826980710e-08 wdrout = -4.026333161e-06 pdrout = 1.825006329e-12
+ pscbe1 = 8.626304063e+08 lpscbe1 = -2.293712868e+01 wpscbe1 = -6.256272284e+03 ppscbe1 = 2.291234098e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 9.095149961e-08 lalpha0 = -2.571138738e-13 walpha0 = -6.088563054e-12 palpha0 = 2.568360159e-17
+ alpha1 = 8.449063844e-01 lalpha1 = 2.601747532e-09 walpha1 = 5.088111020e-07 palpha1 = -2.598935876e-13
+ beta0 = 1.381870533e+01 lbeta0 = -1.658996662e-07 wbeta0 = 4.125004454e-06 pbeta0 = 1.657203817e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.088932651e-01 lkt1 = -9.493876666e-09 wkt1 = 2.780952962e-07 pkt1 = 3.653798084e-14
+ kt2 = -4.863894634e-02 lkt2 = 7.262486249e-10 wkt2 = 2.215918350e-07 pkt2 = -7.397270157e-14
+ at = 1.724245120e+05 lat = -2.703388781e-02 wat = -6.816543185e-01 pat = 1.155914950e-7
+ ute = -2.117471039e+00 lute = 1.947336395e-07 wute = 1.228547208e-05 pute = -5.187023334e-12
+ ua1 = -3.889710299e-10 lua1 = 4.224620078e-16 wua1 = 2.548682287e-14 pua1 = -1.060853673e-20
+ ub1 = -7.957208323e-20 lub1 = -2.241104874e-25 wub1 = -1.145746394e-23 pub1 = 3.455141541e-30
+ uc1 = 1.652876450e-11 luc1 = 1.206696827e-17 wuc1 = 7.610674947e-16 puc1 = -5.783986598e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.6 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.227670599e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.879237320e-09 wvth0 = 7.708900208e-07 pvth0 = -1.877206466e-13
+ k1 = 5.759751139e-01 lk1 = -1.089845111e-08 wk1 = -2.606171909e-06 pk1 = 1.088667337e-12
+ k2 = -4.265052859e-02 lk2 = 3.439071106e-09 wk2 = 8.557384789e-07 pk2 = -3.435354570e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.625148754e-01 ldsub = -6.413663034e-09 wdsub = -2.512157659e-07 pdsub = 6.406731917e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.001421779e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.180212539e-10 wvoff = -1.773543439e-07 pvoff = -3.176775747e-14
+ nfactor = 2.789046350e+00 lnfactor = -1.237454362e-08 wnfactor = -1.815670767e-06 pnfactor = 1.236117070e-12
+ eta0 = -3.577527649e-02 weta0 = 3.623607453e-6
+ etab = -5.592675218e-04 letab = 2.279648880e-11 wetab = 5.851314939e-09 petab = -2.277185309e-15
+ u0 = 2.914241571e-02 lu0 = 3.169428958e-10 wu0 = 2.483156476e-08 pu0 = -3.166003820e-14
+ ua = -9.139636730e-10 lua = 2.032957240e-17 wua = -1.096593353e-15 pua = -2.030760264e-21
+ ub = 1.603607069e-18 lub = -9.841882920e-27 wub = 2.467623486e-24 pub = 9.831246994e-31
+ uc = 7.383107134e-11 luc = -7.261444363e-20 wuc = 4.824067653e-17 puc = 7.253597065e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.068210421e+04 lvsat = -1.926829592e-03 wvsat = -6.813670751e-02 pvsat = 1.924747306e-7
+ a0 = 1.271247476e+00 wa0 = 1.576546842e-6
+ ags = 3.928289067e-01 lags = 4.858609127e-08 wags = 1.475374800e-05 pags = -4.853358525e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.481237729e-04 lketa = 4.622421863e-10 wketa = -1.074281562e-07 pketa = -4.617426504e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.511882494e-01 lpclm = 4.920329430e-09 wpclm = 7.953146481e-07 ppclm = -4.915012128e-13
+ pdiblc1 = 2.766248118e-01 lpdiblc1 = 3.482030347e-08 wpdiblc1 = 1.132526659e-05 ppdiblc1 = -3.478267387e-12
+ pdiblc2 = 4.846842543e-03 lpdiblc2 = 3.496388620e-11 wpdiblc2 = -3.431202270e-09 ppdiblc2 = -3.492610142e-15
+ pdiblcb = -4.046081186e-02 lpdiblcb = 7.897166246e-09 wpdiblcb = 1.544410367e-06 ppdiblcb = -7.888631936e-13
+ drout = 6.032873391e-01 ldrout = -1.979217853e-08 wdrout = -4.324055932e-06 pdrout = 1.977078952e-12
+ pscbe1 = 8.362144241e+08 lpscbe1 = -9.444214796e+00 wpscbe1 = -3.617528787e+03 ppscbe1 = 9.434008622e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.721592095e-07 lalpha0 = 1.326723929e-13 walpha0 = 7.014004001e-11 palpha0 = -1.325290165e-17
+ alpha1 = 0.85
+ beta0 = 1.351919086e+01 lbeta0 = -1.291186681e-08 wbeta0 = 3.404408377e-05 pbeta0 = 1.289791322e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.286328252e-01 lkt1 = 5.888142947e-10 wkt1 = 4.647796970e-07 pkt1 = -5.881779749e-14
+ kt2 = -4.751653897e-02 lkt2 = 1.529386538e-10 wkt2 = 1.066799855e-07 pkt2 = -1.527733760e-14
+ at = 1.173723186e+05 lat = 1.086001837e-03 wat = -2.429690048e-01 pat = -1.084828216e-7
+ ute = -1.693075960e+00 lute = -2.204142494e-08 wute = -2.180045486e-06 pute = 2.201760521e-12
+ ua1 = 4.642273863e-10 lua1 = -1.333979846e-17 wua1 = 2.108979768e-15 pua1 = 1.332538240e-21
+ ub1 = -4.849345502e-19 lub1 = -1.705701435e-26 wub1 = -8.028858962e-24 pub1 = 1.703858118e-30
+ uc1 = 4.817616651e-11 luc1 = -4.098081613e-18 wuc1 = -1.172744218e-15 puc1 = 4.093652898e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.7 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.223204654e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.995702910e-09 wvth0 = 8.155012068e-07 pvth0 = -1.993546193e-13
+ k1 = 5.594265456e-01 lk1 = -6.582816168e-09 wk1 = -9.531034461e-07 pk1 = 6.575702251e-13
+ k2 = -3.909373375e-02 lk2 = 2.511508806e-09 wk2 = 5.004433705e-07 pk2 = -2.508794669e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.058087301e-01 ldsub = 8.374505792e-09 wdsub = 5.413270651e-06 pdsub = -8.365455631e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.014532215e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.599230758e-10 wvoff = -4.639166355e-08 pvoff = -6.592099101e-14
+ nfactor = 2.754218570e+00 lnfactor = -3.291946142e-09 wnfactor = 1.663343481e-06 pnfactor = 3.288388602e-13
+ eta0 = -1.284871776e-01 leta0 = 2.417796585e-08 weta0 = 1.288477838e-05 peta0 = -2.415183720e-12
+ etab = -6.019751828e-03 letab = 1.446814349e-09 wetab = 5.513096419e-07 petab = -1.445250806e-13
+ u0 = 3.359495311e-02 lu0 = -8.442165210e-10 wu0 = -4.199409978e-07 pu0 = 8.433041931e-14
+ ua = -5.614905365e-10 lua = -7.159048698e-17 wua = -3.630581594e-14 pua = 7.151312057e-21
+ ub = 1.389162684e-18 lub = 4.608221042e-26 wub = 2.388888739e-23 pub = -4.603241030e-30
+ uc = 7.391841099e-11 luc = -9.539139970e-20 wuc = 3.951615088e-17 puc = 9.528831212e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.363106444e+04 lvsat = -8.801713357e-05 wvsat = 6.362052782e-01 pvsat = 8.792201522e-9
+ a0 = 1.271247476e+00 wa0 = 1.576546842e-6
+ ags = 8.276643286e-01 lags = -6.481289906e-08 wags = -2.868280239e-05 pags = 6.474285706e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.581967936e-03 lketa = 3.615850247e-11 wketa = -2.706360062e-07 pketa = -3.611942670e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.446950564e-01 lpclm = 6.613663250e-09 wpclm = 1.443932238e-06 ppclm = -6.606515997e-13
+ pdiblc1 = 4.619969338e-01 lpdiblc1 = -1.352215071e-08 wpdiblc1 = -7.191912812e-06 ppdiblc1 = 1.350753760e-12
+ pdiblc2 = 6.251297878e-03 lpdiblc2 = -3.312984028e-10 wpdiblc2 = -1.437249591e-07 ppdiblc2 = 3.309403752e-14
+ pdiblcb = 1.782452985e-02 lpdiblcb = -7.302834878e-09 wpdiblcb = -4.277825024e-06 ppdiblcb = 7.294942850e-13
+ drout = 4.702130150e-01 ldrout = 1.491174215e-08 wdrout = 8.968995400e-06 pdrout = -1.489562733e-12
+ pscbe1 = 7.991711766e+08 lpscbe1 = 2.161455343e-01 wpscbe1 = 8.279276883e+01 ppscbe1 = -2.159119501e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.946638415e-07 lalpha0 = 1.385412859e-13 walpha0 = 7.238807117e-11 palpha0 = -1.383915671e-17
+ alpha1 = 9.188950814e-01 lalpha1 = -1.796687269e-08 walpha1 = -6.882062782e-06 palpha1 = 1.794745625e-12
+ beta0 = 1.263611164e+01 lbeta0 = 2.173828308e-07 wbeta0 = 1.222565732e-04 pbeta0 = -2.171479095e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.198038924e-01 lkt1 = -1.713647765e-09 wkt1 = -4.171594542e-07 pkt1 = 1.711795860e-13
+ kt2 = -4.616455406e-02 lkt2 = -1.996400831e-10 wkt2 = -2.837239922e-08 pkt2 = 1.994243361e-14
+ at = 1.235649369e+05 lat = -5.289463121e-04 wat = -8.615616081e-01 pat = 5.283746904e-8
+ ute = -1.970598865e+00 lute = 5.033266315e-08 wute = 2.554225359e-05 pute = -5.027826965e-12
+ ua1 = 5.995254285e-12 lua1 = 1.061607263e-16 wua1 = 4.788267274e-14 pua1 = -1.060460006e-20
+ ub1 = -2.101392518e-19 lub1 = -8.871978104e-26 wub1 = -3.547869222e-23 pub1 = 8.862390335e-30
+ uc1 = 4.085764812e-11 luc1 = -2.189514478e-18 wuc1 = -4.416832776e-16 puc1 = 2.187148314e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.8 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.268831981e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.125197404e-09 wvth0 = 3.597210303e-07 pvth0 = -1.123981426e-13
+ k1 = 5.312785764e-01 lk1 = -1.212577708e-09 wk1 = 1.858651584e-06 pk1 = 1.211267300e-13
+ k2 = -3.087042946e-02 lk2 = 9.426174735e-10 wk2 = -3.209983826e-07 pk2 = -9.415988056e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.209432474e-01 ldsub = 5.487051776e-09 wdsub = 3.901454479e-06 pdsub = -5.481122029e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 3.255239980e-03 lcdscd = 4.091902473e-10 wcdscd = 2.142442546e-07 pcdscd = -4.087480436e-14
+ cit = 0.0
+ voff = {-1.230164554e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.773886218e-09 wvoff = 2.107601431e-06 pvoff = -4.768727175e-13
+ nfactor = 1.877145382e+00 lnfactor = 1.640413391e-07 wnfactor = 8.927587873e-05 pnfactor = -1.638640629e-11
+ eta0 = -1.375413602e-02 leta0 = 2.288507773e-09 weta0 = 1.423873186e-06 peta0 = -2.286034628e-13
+ etab = -4.088343487e-03 letab = 1.078328677e-09 wetab = 3.583775313e-07 petab = -1.077163349e-13
+ u0 = 2.412533861e-02 lu0 = 9.624533496e-10 wu0 = 5.259970892e-07 pu0 = -9.614132455e-14
+ ua = -1.561762283e-09 lua = 1.192473585e-16 wua = 6.361326137e-14 pua = -1.191184903e-20
+ ub = 2.182599896e-18 lub = -1.052945015e-25 wub = -5.536908863e-23 pub = 1.051807118e-29
+ uc = 6.020391540e-11 luc = 2.521142355e-18 wuc = 1.409483611e-15 puc = -2.518417807e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.953013081e+04 lvsat = -1.213476411e-03 wvsat = 4.693614096e-02 pvsat = 1.212165031e-7
+ a0 = 1.271247476e+00 wa0 = 1.576546842e-6
+ ags = 4.879491552e-01 wags = 5.252002603e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.729722354e-02 lketa = -4.679166254e-09 wketa = -2.739490639e-06 pketa = 4.674109572e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.329144285e-01 lpclm = 8.861242133e-09 wpclm = 2.620721924e-06 ppclm = -8.851665966e-13
+ pdiblc1 = 3.958216889e-01 lpdiblc1 = -8.968404512e-10 wpdiblc1 = -5.815397536e-07 ppdiblc1 = 8.958712537e-14
+ pdiblc2 = 4.801725630e-03 lpdiblc2 = -5.474031191e-11 wpdiblc2 = 1.075613326e-09 ppdiblc2 = 5.468115515e-15
+ pdiblcb = 1.384183335e-02 lpdiblcb = -6.542992142e-09 wpdiblcb = -3.879985776e-06 ppdiblcb = 6.535921262e-13
+ drout = 4.767543002e-01 ldrout = 1.366375651e-08 wdrout = 8.315573786e-06 pdrout = -1.364899037e-12
+ pscbe1 = 7.981748633e+08 lpscbe1 = 4.062281646e-01 wpscbe1 = 1.823164298e+02 ppscbe1 = -4.057891619e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.951900711e-08 lalpha0 = -1.530523077e-15 walpha0 = -9.508720107e-13 palpha0 = 1.528869071e-19
+ alpha1 = 6.892448102e-01 lalpha1 = 2.584718395e-08 walpha1 = 1.605814649e-05 palpha1 = -2.581925142e-12
+ beta0 = 1.332273551e+01 lbeta0 = 8.638460776e-08 wbeta0 = 5.366838757e-05 pbeta0 = -8.629125364e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.114258703e-01 lkt1 = -3.312057091e-09 wkt1 = -1.254056269e-06 pkt1 = 3.308477817e-13
+ kt2 = -4.453891522e-02 lkt2 = -5.097892149e-10 wkt2 = -1.907606037e-07 pkt2 = 5.092382959e-14
+ at = 1.195066423e+05 lat = 2.453194799e-04 wat = -4.561707207e-01 pat = -2.450543680e-8
+ ute = -9.821497330e-01 lute = -1.382495928e-07 wute = -7.319583984e-05 pute = 1.381001893e-11
+ ua1 = 1.571650889e-09 lua1 = -1.925444496e-16 wua1 = -1.085136935e-13 pua1 = 1.923363707e-20
+ ub1 = -1.253525650e-18 lub1 = 1.103437364e-25 wub1 = 6.874719095e-23 pub1 = -1.102244901e-29
+ uc1 = 4.017607318e-11 luc1 = -2.059479521e-18 wuc1 = -3.735994396e-16 puc1 = 2.057253882e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.9 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.188593681e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.772767157e-07 wvth0 = -1.910766174e-08 pvth0 = 1.910972270e-12
+ k1 = 5.418064353e-01 lk1 = -9.408868149e-08 wk1 = -6.483828602e-09 pk1 = 6.484527948e-13
+ k2 = -2.769247282e-02 lk2 = 9.842879788e-08 wk2 = 6.782914213e-09 pk2 = -6.783645819e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.045417318e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.269465504e-08 wvoff = -5.009525865e-09 pvoff = 5.010066193e-13
+ nfactor = 2.550155693e+00 lnfactor = 1.343888008e-05 wnfactor = 9.260985874e-07 pnfactor = -9.261984764e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.149477126e-02 lu0 = -3.267478013e-09 wu0 = -2.251680762e-10 pu0 = 2.251923628e-14
+ ua = -7.366463064e-10 lua = -2.131506240e-15 wua = -1.468861175e-16 pua = 1.469019606e-20
+ ub = 1.537372114e-18 lub = 3.312145784e-24 wub = 2.282462165e-25 pub = -2.282708352e-29
+ uc = 4.773753148e-11 luc = 1.504630793e-16 wuc = 1.036869474e-17 puc = -1.036981311e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.376452071e+00 la0 = -7.001826012e-07 wa0 = -4.825090441e-08 pa0 = 4.825610875e-12
+ ags = 3.811550339e-01 lags = -1.130155785e-07 wags = -7.788116792e-09 pags = 7.788956818e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 8.180254810e-25 lb1 = 1.289455985e-28 wb1 = 8.885884532e-30 pb1 = -8.886842964e-34
+ keta = -7.199184736e-03 lketa = -1.595587346e-07 wketa = -1.099549351e-08 pketa = 1.099667949e-12
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.725335471e-02 lpclm = -3.094069161e-06 wpclm = -2.132181449e-07 ppclm = 2.132411426e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.147018095e-03 lpdiblc2 = -7.356732866e-09 wpdiblc2 = -5.069663451e-10 ppdiblc2 = 5.070210265e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.178768667e+08 lpscbe1 = 3.680126221e+03 wpscbe1 = 2.536044429e+02 ppscbe1 = -2.536317966e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.199864079e-01 lkt1 = 6.957158242e-07 wkt1 = 4.794309037e-08 pkt1 = -4.794826152e-12
+ kt2 = -4.543335553e-02 lkt2 = 1.200314779e-08 wkt2 = 8.271595661e-10 pkt2 = -8.272487835e-14
+ at = 140000.0
+ ute = -1.856411036e+00 lute = 4.301567497e-06 wute = 2.964291340e-07 pute = -2.964611068e-11
+ ua1 = 3.044858563e-10 lua1 = 7.154185942e-15 wua1 = 4.930084544e-16 pua1 = -4.930616303e-20
+ ub1 = -5.528820975e-19 lub1 = -8.674725804e-24 wub1 = -5.977917258e-25 pub1 = 5.978562036e-29
+ uc1 = 1.656219400e-11 luc1 = -7.325600042e-17 wuc1 = -5.048209235e-18 puc1 = 5.048753735e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.10 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.050030051e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 7.638945015e-8
+ k1 = 5.371045370e-01 wk1 = 2.592133503e-8
+ k2 = -2.277368563e-02 wk2 = -2.711703264e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.081745054e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 2.002730274e-8
+ nfactor = 3.221737513e+00 wnfactor = -3.702397647e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.133148542e-02 wu0 = 9.001868339e-10
+ ua = -8.431641733e-10 wua = 5.872277781e-16
+ ub = 1.702890140e-18 wub = -9.124927588e-25
+ uc = 5.525663039e-11 wuc = -4.145242368e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.341461811e+00 wa0 = 1.928995869e-7
+ ags = 3.755073008e-01 wags = 3.113567570e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 7.261830261e-24 wb1 = -3.552437983e-29
+ keta = -1.517282128e-02 wketa = 4.395826736e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.736671676e-02 wpclm = 8.524128735e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.779379719e-03 wpdiblc2 = 2.026772342e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 9.017839967e+08 wpscbe1 = -1.013870991e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.852193666e-01 wkt1 = -1.916689944e-7
+ kt2 = -4.483352163e-02 wkt2 = -3.306854877e-9
+ at = 140000.0
+ ute = -1.641448590e+00 wute = -1.185077424e-6
+ ua1 = 6.620023447e-10 wua1 = -1.970970873e-15
+ ub1 = -9.863845998e-19 wub1 = 2.389878042e-24
+ uc1 = 1.290136826e-11 wuc1 = 2.018195281e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.11 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.865892412e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.475087222e-07 wvth0 = 1.471195825e-07 pvth0 = -5.666039541e-13
+ k1 = 5.246957231e-01 lk1 = 9.940435247e-08 wk1 = 4.822739943e-08 pk1 = -1.786891084e-13
+ k2 = -1.122526934e-02 lk2 = -9.251189154e-08 wk2 = -6.859979467e-08 pk2 = 3.323095293e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.176113977e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.559692437e-08 wvoff = 6.005283304e-08 pvoff = -3.206359578e-13
+ nfactor = 3.787202708e+00 lnfactor = -4.529820674e-06 wnfactor = -7.739483276e-06 pnfactor = 3.234022904e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.189532637e-02 lu0 = -4.516809250e-09 wu0 = 6.263600579e-10 pu0 = 2.193567704e-15
+ ua = -8.804820293e-10 lua = 2.989453581e-16 wua = 8.064207034e-16 pua = -1.755907617e-21
+ ub = 1.877153765e-18 lub = -1.395988610e-24 wub = -1.585058649e-24 pub = 5.387781416e-30
+ uc = 1.749290886e-10 luc = -9.586704525e-16 wuc = -8.223658220e-16 puc = 6.255730119e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.769452386e+00 la0 = -3.428540902e-06 wa0 = -2.039645614e-06 pa0 = 1.788444184e-11
+ ags = 4.476107193e-01 lags = -5.776050552e-07 wags = -6.188986654e-07 pags = 5.207285999e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 1.454324205e-23 lb1 = -5.832983160e-29 wb1 = -7.114455115e-29 pb1 = 2.853455697e-34
+ keta = -2.844591055e-02 lketa = 1.063278777e-07 wketa = 8.835622306e-08 pketa = -3.556625219e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.020884212e+00 lpclm = 7.398101022e-06 wpclm = 3.342478635e-06 ppclm = -1.994738394e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 2.818096188e-03 lpdiblc2 = -3.101493542e-10 wpdiblc2 = 1.641582583e-09 ppdiblc2 = 3.085672732e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.001221352e+09 lpscbe1 = -7.965713764e+02 wpscbe1 = -2.012411431e+03 ppscbe1 = 7.999093778e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.601231753e-01 lkt1 = -2.010402180e-07 wkt1 = -3.500490494e-07 pkt1 = 1.268748728e-12
+ kt2 = -3.219755090e-02 lkt2 = -1.012240574e-07 wkt2 = -8.264351494e-08 pkt2 = 6.355490057e-13
+ at = 140000.0
+ ute = -1.123537024e+00 lute = -4.148878724e-06 wute = -4.479450180e-06 pute = 2.639051515e-11
+ ua1 = 1.912795055e-09 lua1 = -1.001983273e-14 wua1 = -9.230253929e-15 pua1 = 5.815256307e-20
+ ub1 = -2.186713527e-18 lub1 = 9.615578161e-24 wub1 = 8.880586807e-24 pub1 = -5.199567891e-29
+ uc1 = -2.771450635e-11 luc1 = 3.253650797e-16 wuc1 = 1.997098526e-16 puc1 = -1.438159586e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.12 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.238910272e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.100759086e-09 wvth0 = -4.119398830e-08 pvth0 = 1.886814793e-13
+ k1 = 5.756552523e-01 lk1 = -1.049834137e-07 wk1 = -1.758356650e-07 pk1 = 7.199798934e-13
+ k2 = -4.225743877e-02 lk2 = 3.195149914e-08 wk2 = 8.205363029e-08 pk2 = -2.719291184e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.871247706e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.031046194e-08 wvoff = -8.729703218e-08 pvoff = 2.703528187e-13
+ nfactor = 2.520055606e+00 lnfactor = 5.524351856e-07 wnfactor = 8.151637335e-07 pnfactor = -1.970629421e-12
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398724195e-01 letab = 2.802433220e-07 wetab = -1.171062741e-11 petab = 4.696882045e-17
+ u0 = 3.207753642e-02 lu0 = -5.247614758e-09 wu0 = 2.885059913e-09 pu0 = -6.865594051e-15
+ ua = -4.011086334e-10 lua = -1.623718747e-15 wua = -1.226352763e-15 pua = 6.397111744e-21
+ ub = 9.744011767e-19 lub = 2.224758832e-24 wub = 2.650668732e-24 pub = -1.160081466e-29
+ uc = -2.093422232e-10 luc = 5.825595450e-16 wuc = 1.520696392e-15 puc = -3.141791005e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 4.153275676e-01 la0 = 2.002563960e-06 wa0 = 5.712583713e-06 pa0 = -1.320809101e-11
+ ags = 1.144642986e-01 lags = 7.585739446e-07 wags = 1.024303754e-06 pags = -1.383247261e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.180386289e-05 lketa = -7.635023608e-09 wketa = -2.629050060e-08 pketa = 1.041609523e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.320634398e-01 lpclm = -3.367547891e-08 wpclm = -1.495708702e-06 ppclm = -5.424499062e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 1.305949366e-03 lpdiblc2 = 5.754747951e-09 wpdiblc2 = 3.683254340e-10 ppdiblc2 = 8.192434679e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.052422032e+08 lpscbe1 = -1.054094871e+01 wpscbe1 = -3.612890767e+01 ppscbe1 = 7.264750173e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.046064812e-01 lkt1 = -2.262719718e-08 wkt1 = -1.134304931e-08 pkt1 = -8.972855592e-14
+ kt2 = -5.800521569e-02 lkt2 = 2.284963183e-09 wkt2 = 7.983863007e-08 pkt2 = -1.613210674e-14
+ at = 1.682199118e+05 lat = -1.131840272e-01 wat = -2.084646247e-02 pat = 8.361069983e-8
+ ute = -2.533092297e+00 lute = 1.504545829e-06 wute = 3.727476919e-06 pute = -6.525713158e-12
+ ua1 = -1.720323789e-09 lua1 = 4.551829464e-15 wua1 = 1.096817911e-14 pua1 = -2.285902938e-20
+ ub1 = 1.238884608e-18 lub1 = -4.123762879e-24 wub1 = -9.897674307e-24 pub1 = 2.331990787e-29
+ uc1 = 6.694697625e-11 luc1 = -5.430186945e-17 wuc1 = -2.942920936e-16 puc1 = 5.431765036e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.13 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.943497501e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.730042734e-08 wvth0 = 7.171955536e-08 pvth0 = -3.836349352e-14
+ k1 = 4.320314661e-01 lk1 = 1.838132848e-07 wk1 = 5.771236946e-07 pk1 = -7.940602453e-13
+ k2 = 1.043823076e-02 lk2 = -7.400821541e-08 wk2 = -2.113560778e-07 pk2 = 3.180550150e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.152362433e+00 ldsub = -1.794349887e-06 wdsub = -6.150101207e-06 pdsub = 1.236653740e-11
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.036330347e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.030841350e-08 wvoff = 1.422205481e-07 pvoff = -1.911579184e-13
+ nfactor = 2.908375480e+00 lnfactor = -2.283929821e-07 wnfactor = -1.331454003e-07 pnfactor = -6.378269137e-14
+ eta0 = -6.590106194e-03 leta0 = 1.425668627e-08 weta0 = 3.471429712e-08 peta0 = -6.980302264e-14
+ etab = -9.758147600e-04 letab = 9.519737058e-10 wetab = 1.963530663e-09 petab = -3.924818713e-15
+ u0 = 3.309312078e-02 lu0 = -7.289737565e-09 wu0 = -7.636131088e-10 pu0 = 4.711065784e-16
+ ua = -9.099793181e-10 lua = -6.004886983e-16 wua = 3.509173667e-15 pua = -3.125018505e-21
+ ub = 1.950124731e-18 lub = 2.627875688e-25 wub = -5.890541933e-24 pub = 5.573732167e-30
+ uc = 7.457786857e-11 luc = 1.165699933e-17 wuc = 9.181504903e-17 puc = -2.686164054e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.885541875e+04 lvsat = 1.229486679e-01 wvsat = 2.799890480e-01 pvsat = -5.629980579e-7
+ a0 = 2.455556164e+00 la0 = -2.099899139e-06 wa0 = -6.731274788e-06 pa0 = 1.181384545e-11
+ ags = 9.420035339e-01 lags = -9.054303641e-07 wags = -5.170032837e-06 pags = 1.107223804e-11
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.356607466e-02 lketa = -1.154088874e-07 wketa = 8.236954313e-08 pketa = -1.143311424e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.101756931e+00 lpclm = -5.759713759e-07 wpclm = -2.572969108e-06 ppclm = 1.623690236e-12
+ pdiblc1 = -2.053601678e-01 lpdiblc1 = 1.197141890e-06 wpdiblc1 = 1.893742697e-06 ppdiblc1 = -3.807911303e-12
+ pdiblc2 = 6.892558304e-03 lpdiblc2 = -5.478727089e-09 wpdiblc2 = -8.755152680e-09 ppdiblc2 = 2.653779674e-14
+ pdiblcb = -4.984180035e-02 lpdiblcb = 4.995154436e-08 wpdiblcb = -1.614028203e-09 ppdiblcb = 3.245465313e-15
+ drout = 8.632358000e-01 ldrout = -6.097423013e-7
+ pscbe1 = 2.367661598e+09 lpscbe1 = -3.152231995e+03 wpscbe1 = -7.049917884e+03 ppscbe1 = 1.417587618e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.586663671e-07 lalpha0 = -6.608777297e-13 walpha0 = -2.044710672e-11 palpha0 = 4.111475594e-17
+ alpha1 = 8.156332760e-01 lalpha1 = 6.910412749e-8
+ beta0 = 1.174294166e+01 lbeta0 = 4.256951278e-06 wbeta0 = -4.719873801e-06 pbeta0 = 9.490656162e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.617030336e-01 lkt1 = 9.218175103e-08 wkt1 = -9.731532246e-08 pkt1 = 8.314328732e-14
+ kt2 = -8.777548880e-02 lkt2 = 6.214661158e-08 wkt2 = 1.450663766e-07 pkt2 = -1.472911463e-13
+ at = 1.579085934e+05 lat = -9.245017255e-02 wat = 6.314170135e-02 pat = -8.527152414e-8
+ ute = -2.589035663e+00 lute = 1.617035967e-06 wute = 2.558505937e-07 pute = 4.549844548e-13
+ ua1 = -9.103542364e-10 lua1 = 2.923154027e-15 wua1 = -2.355051396e-15 pua1 = 3.931135995e-21
+ ub1 = -3.210116898e-19 lub1 = -9.871452416e-25 wub1 = 4.602988815e-24 pub1 = -5.837822523e-30
+ uc1 = 1.085175074e-11 luc1 = 5.849362467e-17 wuc1 = 4.096213043e-17 puc1 = -1.309479965e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.14 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.324359490e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.880343073e-08 wvth0 = -4.246350278e-08 pvth0 = 7.705114309e-14
+ k1 = 7.243968413e-01 lk1 = -1.117055434e-07 wk1 = -2.808983443e-07 pk1 = 7.321641923e-14
+ k2 = -1.117546243e-01 lk2 = 4.950261180e-08 wk2 = 1.701099009e-07 pk2 = -6.752545577e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.760407772e+00 ldsub = 1.149837457e-06 wdsub = 1.297050040e-05 pdsub = -6.960299009e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.065630528e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.346792241e-09 wvoff = -9.486017314e-10 pvoff = -4.644454612e-14
+ nfactor = 2.268773401e+00 lnfactor = 4.181078448e-07 wnfactor = 1.256550378e-06 pnfactor = -1.468467728e-12
+ eta0 = -4.853792816e-01 leta0 = 4.982100817e-07 weta0 = -6.942859423e-08 peta0 = 3.546315393e-14
+ etab = 2.505088655e-04 letab = -2.875770464e-10 wetab = -3.880218816e-09 petab = 1.981961448e-15
+ u0 = 2.852315666e-02 lu0 = -2.670481817e-09 wu0 = -8.186854767e-09 pu0 = 7.974415321e-15
+ ua = -1.260373075e-09 lua = -2.463155942e-16 wua = -8.855258609e-17 pua = 5.115128236e-22
+ ub = 2.114752812e-18 lub = 9.638380952e-26 wub = -1.848191152e-25 pub = -1.935325775e-31
+ uc = 8.651100948e-11 luc = -4.048524357e-19 wuc = -3.307156876e-16 puc = 1.584717478e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.818236357e+05 lvsat = -4.177732423e-02 wvsat = -7.125172551e-01 pvsat = 4.402134182e-7
+ a0 = -7.680726914e-01 la0 = 1.158499778e-06 wa0 = 1.001993426e-05 pa0 = -5.118042139e-12
+ ags = -1.183497760e+00 lags = 1.242996587e-06 wags = 1.169288245e-05 pags = -5.972560655e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.287715622e-02 lketa = 2.250602020e-08 wketa = -1.463844231e-07 pketa = 1.168901641e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.454808005e-01 lpclm = 2.895405492e-07 wpclm = -1.272950021e-08 ppclm = -9.641641155e-13
+ pdiblc1 = 6.539326663e-01 lpdiblc1 = 3.285807237e-07 wpdiblc1 = -1.694896701e-06 ppdiblc1 = -1.805648400e-13
+ pdiblc2 = -1.581019058e-03 lpdiblc2 = 3.086246279e-09 wpdiblc2 = 4.266929097e-08 ppdiblc2 = -2.544131096e-14
+ pdiblcb = 2.468360070e-02 lpdiblcb = -2.537768767e-08 wpdiblcb = 3.228056405e-09 ppdiblcb = -1.648846019e-15
+ drout = 1.061865782e+00 ldrout = -8.105147058e-07 wdrout = -7.207365652e-06 pdrout = 7.285104298e-12
+ pscbe1 = -1.493337837e+09 lpscbe1 = 7.504121807e+02 wpscbe1 = 9.980900644e+03 ppscbe1 = -3.038636754e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.164353793e-05 lalpha0 = 2.157864235e-11 walpha0 = 1.437040602e-10 palpha0 = -1.248069455e-16
+ alpha1 = 9.187334480e-01 lalpha1 = -3.510808297e-8
+ beta0 = 7.038229371e-01 lbeta0 = 1.541513793e-05 wbeta0 = 9.451188209e-05 pbeta0 = -9.081141345e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.685231124e-01 lkt1 = -2.003208800e-09 wkt1 = -1.330503908e-10 pkt1 = -1.508719273e-14
+ kt2 = -1.693659162e-02 lkt2 = -9.456353950e-09 wkt2 = 3.101362028e-09 pkt2 = -3.794897042e-15
+ at = 8.077706654e+04 lat = -1.448670502e-02 wat = -5.002635658e-02 pat = 2.911716446e-8
+ ute = -6.535547181e-01 lute = -3.393210752e-07 wute = 2.196260345e-06 pute = -1.506354556e-12
+ ua1 = 2.635044555e-09 lua1 = -6.604854357e-16 wua1 = 4.645513098e-15 pua1 = -3.144936588e-21
+ ub1 = -1.241995230e-18 lub1 = -5.622797294e-26 wub1 = -3.446122658e-24 pub1 = 2.298106667e-30
+ uc1 = 1.553485586e-10 luc1 = -8.756172578e-17 wuc1 = -1.956690866e-16 puc1 = 1.082355248e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.15 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.200995669e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.597391799e-08 wvth0 = 1.000810017e-07 pvth0 = 4.241405832e-15
+ k1 = 2.473628332e-01 lk1 = 1.319567495e-07 wk1 = -3.413984157e-07 pk1 = 1.041190087e-13
+ k2 = 6.991576078e-02 lk2 = -4.329207752e-08 wk2 = 7.993926712e-08 pk2 = -2.146755842e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.694105324e-01 ldsub = 6.195608480e-08 wdsub = -9.879333645e-07 pdsub = 1.694735387e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.007302728e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.032609460e-08 wvoff = -1.733012334e-07 pvoff = 4.159076517e-14
+ nfactor = 2.938532925e+00 lnfactor = 7.600405702e-08 wnfactor = -2.845922071e-06 pnfactor = 6.270177640e-13
+ eta0 = 0.49
+ etab = -2.414997841e-04 letab = -3.626591627e-11 wetab = 3.661281299e-09 petab = -1.870131230e-15
+ u0 = 2.953985264e-02 lu0 = -3.189795891e-09 wu0 = 2.209245645e-08 pu0 = -7.491832939e-15
+ ua = -1.304151342e-09 lua = -2.239542685e-16 wua = 1.592553528e-15 pua = -3.471726437e-22
+ ub = 1.901068449e-18 lub = 2.055307907e-25 wub = 4.175398844e-25 pub = -5.012091215e-31
+ uc = -7.331682434e-12 luc = 4.752868080e-17 wuc = 6.076088565e-16 puc = -3.208112929e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.168760594e+04 lvsat = 4.512577789e-02 wvsat = 4.073686830e-01 pvsat = -1.318086406e-7
+ a0 = 1.5
+ ags = 2.533556992e+00 lags = -6.556229419e-07 wags = -4.396182092e-12 pags = 2.245508265e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.321862732e-02 lketa = -7.966721141e-09 wketa = 5.912744897e-08 pketa = 1.191757704e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.264088925e+00 lpclm = -2.307502202e-07 wpclm = -4.117948330e-06 ppclm = 1.132724189e-12
+ pdiblc1 = 3.500271335e+00 lpdiblc1 = -1.125289220e-06 wpdiblc1 = -1.089188604e-05 ppdiblc1 = 4.517128559e-12
+ pdiblc2 = 6.445527389e-03 lpdiblc2 = -1.013601275e-09 wpdiblc2 = -1.444922952e-08 ppdiblc2 = 3.734029647e-15
+ pdiblcb = 6.939277514e-01 lpdiblcb = -3.672182304e-07 wpdiblcb = -3.516945673e-06 ppdiblcb = 1.796406612e-12
+ drout = -2.115658123e+00 ldrout = 8.125200193e-07 wdrout = 1.441473130e-05 pdrout = -3.759160118e-12
+ pscbe1 = -8.839707193e+08 lpscbe1 = 4.391559880e+02 wpscbe1 = 8.237870249e+03 ppscbe1 = -2.148321231e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 4.408558481e-05 lalpha0 = -1.199487334e-11 walpha0 = -2.383272882e-10 palpha0 = 7.032931888e-17
+ alpha1 = 0.85
+ beta0 = 4.385311210e+01 lbeta0 = -6.624914882e-06 wbeta0 = -1.750152387e-04 pbeta0 = 4.685926649e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.062179859e-01 lkt1 = -3.382779518e-08 wkt1 = -3.788950514e-07 pkt1 = 1.783791347e-13
+ kt2 = 3.728318971e-03 lkt2 = -2.001170097e-08 wkt2 = -2.464960908e-07 pkt2 = 1.236959875e-13
+ at = 8.326673287e+04 lat = -1.575839172e-02 wat = -7.915627080e-03 pat = 7.607593381e-9
+ ute = -1.207134136e+00 lute = -5.656045848e-08 wute = -5.529123494e-06 pute = 2.439663353e-12
+ ua1 = 1.794695167e-09 lua1 = -2.312467333e-16 wua1 = -7.060513702e-15 pua1 = 2.834338018e-21
+ ub1 = -2.211127900e-18 lub1 = 4.387914272e-25 wub1 = 3.867948226e-24 pub1 = -1.437818344e-30
+ uc1 = -1.537784305e-10 luc1 = 7.033601246e-17 wuc1 = 2.191131311e-16 puc1 = -1.036294250e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.16 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.773691330e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.483041907e-08 wvth0 = 4.361095333e-07 pvth0 = -8.339013080e-14
+ k1 = 3.929471458e-01 lk1 = 9.399039896e-08 wk1 = 1.942612567e-07 pk1 = -3.557353461e-14
+ k2 = 5.258147608e-02 lk2 = -3.877153875e-08 wk2 = -1.313759417e-07 pk2 = 3.364048963e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.149386476e+00 ldsub = -1.414507217e-07 wdsub = -1.089803013e-06 pdsub = 1.960397170e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-4.391585505e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.514249935e-08 wvoff = -4.429352804e-07 pvoff = 1.119075498e-13
+ nfactor = 4.317577045e+00 lnfactor = -2.836313430e-07 wnfactor = -9.111216819e-06 pnfactor = 2.260918920e-12
+ eta0 = 1.785091854e+00 leta0 = -3.377418242e-07 weta0 = -3.034781852e-07 peta0 = 7.914286201e-14
+ etab = 9.694732365e-02 letab = -2.538175042e-08 wetab = -1.583324405e-07 petab = 4.037556351e-14
+ u0 = -3.158093251e-02 lu0 = 1.274964919e-08 wu0 = 2.924677390e-08 pu0 = -9.357578770e-15
+ ua = -5.801454442e-09 lua = 9.488794177e-16 wua = -1.923410210e-16 pua = 1.183028660e-22
+ ub = 4.365278260e-18 lub = -4.371006291e-25 wub = 3.377701223e-24 pub = -1.273177756e-30
+ uc = 3.824859231e-10 luc = -5.413029328e-17 wuc = -2.087110160e-15 puc = 3.819337006e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.305653097e+05 lvsat = 1.412413704e-02 wvsat = 2.438183315e-01 pvsat = -8.915699862e-8
+ a0 = 1.5
+ ags = -3.334132116e+00 lags = 8.745882298e-07 wags = 1.570065032e-11 pags = -2.995464273e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.252174902e-01 lketa = 1.863315431e-08 wketa = 6.101491687e-07 pketa = -1.317811732e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.344731062e+00 lpclm = -2.517805605e-07 wpclm = -4.069861508e-06 ppclm = 1.120183820e-12
+ pdiblc1 = -4.053430367e+00 lpdiblc1 = 8.446104324e-07 wpdiblc1 = 2.392810509e-05 ppdiblc1 = -4.563437650e-12
+ pdiblc2 = -1.144466001e-02 lpdiblc2 = 3.651909135e-09 wpdiblc2 = -2.176562067e-08 ppdiblc2 = 5.642042029e-15
+ pdiblcb = -2.557604613e+00 lpdiblcb = 4.807358888e-07 wpdiblcb = 1.347185750e-05 ppdiblcb = -2.634035412e-12
+ drout = 2.345302393e+00 ldrout = -3.508360297e-07 wdrout = -3.953993084e-06 pdrout = 1.031146040e-12
+ pscbe1 = 8.224207200e+08 lpscbe1 = -5.847009874e+00 wpscbe1 = -7.744150286e+01 ppscbe1 = 2.019565977e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 4.292487415e-06 lalpha0 = -1.617390645e-12 walpha0 = 3.801696384e-11 palpha0 = -1.737393242e-18
+ alpha1 = -3.544460907e+00 lalpha1 = 1.146013882e-06 walpha1 = 2.387908318e-05 palpha1 = -6.227330586e-12
+ beta0 = 5.046385996e+01 lbeta0 = -8.348905373e-06 wbeta0 = -1.384496959e-04 pbeta0 = 3.732348484e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.365837245e-01 lkt1 = 7.840556432e-08 wkt1 = 1.766065607e-06 pkt1 = -3.809965756e-13
+ kt2 = -1.719377854e-01 lkt2 = 2.579955974e-08 wkt2 = 8.384481588e-07 pkt2 = -1.592422836e-13
+ at = 4.137853949e+04 lat = -4.834537323e-03 wat = -2.951385460e-01 pat = 8.251130951e-8
+ ute = -3.947397095e-01 lute = -2.684215515e-07 wute = 1.468153945e-05 pute = -2.830994593e-12
+ ua1 = 4.987087401e-09 lua1 = -1.063777934e-15 wua1 = 1.355332439e-14 pua1 = -2.541462362e-21
+ ub1 = -5.369234270e-18 lub1 = 1.262381355e-24 wub1 = 7.743982681e-26 pub1 = -4.493068204e-31
+ uc1 = -1.445876184e-10 luc1 = 6.793917735e-17 wuc1 = 8.363928891e-16 puc1 = -2.646073440e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.17 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.090196161e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.790288133e-09 wvth0 = 4.828356227e-07 pvth0 = -9.230481450e-14
+ k1 = 7.799027841e-01 lk1 = 2.016468055e-08 wk1 = 1.451504503e-07 pk1 = -2.620388030e-14
+ k2 = 2.244796591e-03 lk2 = -2.916800502e-08 wk2 = -5.492262687e-07 pk2 = 1.133604821e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.710797545e+00 ldsub = -2.485600938e-07 wdsub = -6.366520028e-06 pdsub = 1.202763449e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 7.964700865e-02 lcdscd = -1.416528827e-08 wcdscd = -3.122425678e-07 pcdscd = 5.957151054e-14
+ cit = 0.0
+ voff = {7.479338327e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.762163339e-07 wvoff = -3.894928730e-06 pvoff = 7.704995720e-13
+ nfactor = 3.897148618e+01 lnfactor = -6.895112052e-06 wnfactor = -1.663757957e-04 pnfactor = 3.226479886e-11
+ eta0 = 8.920538562e-02 leta0 = -1.419042847e-08 weta0 = 7.142831643e-07 peta0 = -1.150317548e-13
+ etab = 5.455232265e-02 letab = -1.729337776e-08 wetab = -4.576995217e-08 petab = 1.890021661e-14
+ u0 = 8.506183898e-02 lu0 = -9.504158615e-09 wu0 = 1.060268723e-07 pu0 = -2.400614662e-14
+ ua = 6.472343722e-09 lua = -1.392789439e-15 wua = 8.242749106e-15 pua = -1.490994239e-21
+ ub = -5.052985640e-18 lub = 1.359772267e-24 wub = -5.501925139e-24 pub = 4.209306387e-31
+ uc = 1.931550608e-10 luc = -1.800861539e-17 wuc = 4.931933579e-16 puc = -1.103520864e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.603722756e+05 lvsat = -2.971981476e-02 wvsat = -1.888608824e+00 pvsat = 3.176802486e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.364558697e+00 lketa = 2.550821058e-07 wketa = 6.853085721e-06 pketa = -1.322846066e-12
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.090050787e+00 lpclm = 2.127417293e-07 wpclm = 1.380608783e-05 ppclm = -2.290297050e-12
+ pdiblc1 = -2.583725971e-01 lpdiblc1 = 1.205665408e-07 wpdiblc1 = 3.927122780e-06 ppdiblc1 = -7.475302386e-13
+ pdiblc2 = -1.070763525e-02 lpdiblc2 = 3.511295130e-09 wpdiblc2 = 1.079650739e-07 ppdiblc2 = -1.910875826e-14
+ pdiblcb = -7.100674871e-01 lpdiblcb = 1.282516707e-07 wpdiblcb = 1.109148035e-06 ppdiblcb = -2.754035238e-13
+ drout = -4.276558212e-01 ldrout = 1.782055760e-07 wdrout = 1.454870684e-05 pdrout = -2.498910068e-12
+ pscbe1 = 8.206498117e+08 lpscbe1 = -5.509145379e+00 wpscbe1 = 2.742061355e+01 ppscbe1 = 1.894360245e-7
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.677559070e-05 lalpha0 = 4.309963707e-12 walpha0 = 1.838570407e-10 palpha0 = -2.956163814e-17
+ alpha1 = 1.110374212e+01 lalpha1 = -1.648658180e-06 walpha1 = -5.571786075e-05 palpha1 = 8.958651959e-12
+ beta0 = -3.165337823e+01 lbeta0 = 7.317914033e-06 wbeta0 = 3.636407051e-04 pbeta0 = -5.846833442e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.083167237e-01 lkt1 = 7.301261631e-08 wkt1 = 7.920953037e-07 pkt1 = -1.951766773e-13
+ kt2 = -7.241605716e-02 lkt2 = 6.812207284e-09 wkt2 = 1.366762845e-09 pkt2 = 4.611276186e-16
+ at = 2.684615213e+05 lat = -4.815879108e-02 wat = -1.482757618e+00 pat = 3.090924017e-7
+ ute = -1.145774539e+01 lute = 1.842245050e-06 wute = -9.987469154e-07 pute = 1.605845215e-13
+ ua1 = -1.664587276e-08 lua1 = 3.063488002e-15 wua1 = 1.704024069e-14 pua1 = -3.206717175e-21
+ ub1 = 9.878810420e-18 lub1 = -1.646732099e-24 wub1 = -7.976112251e-24 pub1 = 1.087198166e-30
+ uc1 = 2.491233437e-10 luc1 = -7.175362263e-18 wuc1 = -1.813649820e-15 puc1 = 2.409837042e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.18 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.156258977e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.610520623e-08 wvth0 = -3.289744144e-09 pvth0 = 3.290098976e-13
+ k1 = 5.437593776e-01 lk1 = -2.894039739e-07 wk1 = -1.603748943e-08 pk1 = 1.603921924e-12
+ k2 = -2.747501919e-02 lk2 = 7.668108845e-08 wk2 = 5.719145794e-09 pk2 = -5.719762661e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.061689583e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 9.004554036e-08 wvoff = 2.950755234e-09 pvoff = -2.951073503e-13
+ nfactor = 2.730804721e+00 lnfactor = -4.627971227e-06 wnfactor = 4.237582545e-08 pnfactor = -4.238039611e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.128149898e-02 lu0 = 1.806204949e-08 wu0 = 8.181453732e-10 pu0 = -8.182336184e-14
+ ua = -7.603977722e-10 lua = 2.438965274e-16 wua = -3.069556171e-17 pua = 3.069887253e-21
+ ub = 1.561449713e-18 lub = 9.041262229e-25 wub = 1.104602415e-25 pub = -1.104721557e-29
+ uc = 5.860591513e-11 luc = -9.364925123e-16 wuc = -4.279869903e-17 puc = 4.280331530e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.389986204e+00 la0 = -2.053741873e-06 wa0 = -1.144589624e-07 pa0 = 1.144713079e-11
+ ags = 3.837046725e-01 lags = -3.680069434e-07 wags = -2.026077567e-08 pags = 2.026296099e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.621818611e-25 lb0 = -7.622640700e-29 wb0 = -3.728541836e-30 pb0 = 3.728943997e-34
+ b1 = 2.634462122e-24 lb1 = -5.271765776e-29
+ keta = -9.255513369e-03 lketa = 4.609630834e-08 wketa = -9.360736683e-10 pketa = 9.361746332e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.607253566e-02 lpclm = 1.024456920e-06 wpclm = -1.176437843e-08 ppclm = 1.176564734e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.778937312e-03 lpdiblc2 = 2.945531555e-08 wpdiblc2 = 1.293659815e-09 ppdiblc2 = -1.293799350e-13
+ pdiblcb = -9.243755364e-01 lpdiblcb = 8.994725431e-05 wpdiblcb = 4.399683967e-06 ppdiblcb = -4.400158517e-10
+ drout = 0.56
+ pscbe1 = 8.055199410e+08 lpscbe1 = -5.085126522e+03 wpscbe1 = -1.751395166e+02 ppscbe1 = 1.751584072e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.072707742e-01 lkt1 = -5.759846956e-07 wkt1 = -1.426092497e-08 pkt1 = 1.426246316e-12
+ kt2 = -4.365554522e-02 lkt2 = -1.657970589e-07 wkt2 = -7.869767593e-09 pkt2 = 7.870616426e-13
+ at = 140000.0
+ ute = -1.762034007e+00 lute = -5.137153318e-06 wute = -1.652568725e-07 pute = 1.652746971e-11
+ ua1 = 4.312276173e-10 lua1 = -5.521357198e-15 wua1 = -1.270036222e-16 pua1 = 1.270173208e-20
+ ub1 = -6.487906259e-19 lub1 = 9.171615061e-25 wub1 = -1.286137266e-25 pub1 = 1.286275989e-29
+ uc1 = 1.485765777e-11 luc1 = 9.721600786e-17 wuc1 = 3.290266101e-18 puc1 = -3.290620990e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.19 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.179299154e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.315188377e-8
+ k1 = 5.292969785e-01 wk1 = 6.411538031e-8
+ k2 = -2.364303135e-02 wk2 = -2.286425249e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016691080e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -1.179665900e-8
+ nfactor = 2.499530886e+00 wnfactor = -1.694119379e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.218411468e-02 wu0 = -3.270817541e-9
+ ua = -7.482095190e-10 wua = 1.227160661e-16
+ ub = 1.606631657e-18 wub = -4.416028094e-25
+ uc = 1.180652843e-11 wuc = 1.711025205e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.287354459e+00 wa0 = 4.575890716e-7
+ ags = 3.653142433e-01 wags = 8.099941968e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -3.047084152e-24 wb0 = 1.490612847e-29
+ b1 = 0.0
+ keta = -6.951940269e-03 wketa = 3.742276463e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.726777207e-02 wpclm = 4.703214929e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 4.250909254e-03 wpdiblc2 = -5.171850083e-9
+ pdiblcb = 3.570563059e+00 wpdiblcb = -1.758924998e-5
+ drout = 0.56
+ pscbe1 = 5.514006614e+08 wpscbe1 = 7.001804591e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.360544860e-01 wkt1 = 5.701295281e-8
+ kt2 = -5.194092986e-02 wkt2 = 3.146210286e-8
+ at = 140000.0
+ ute = -2.018753224e+00 wute = 6.606711901e-7
+ ua1 = 1.553085605e-10 wua1 = 5.077406641e-16
+ ub1 = -6.029572685e-19 wub1 = 5.141776104e-25
+ uc1 = 1.971583814e-11 wuc1 = -1.315397047e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.20 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.261220831e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.562570242e-08 wvth0 = -4.627239217e-08 pvth0 = 4.760351578e-13
+ k1 = 5.146731750e-01 lk1 = 1.171481599e-07 wk1 = 9.725702309e-08 pk1 = -2.654906080e-13
+ k2 = -2.136305342e-02 lk2 = -1.826441535e-08 wk2 = -1.900644435e-08 pk2 = -3.090407540e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017764992e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 8.602876988e-10 wvoff = -1.741041360e-08 pvoff = 4.497058676e-14
+ nfactor = 1.645326577e+00 lnfactor = 6.842847914e-06 wnfactor = 2.738429110e-06 pnfactor = -2.329409235e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.350013523e-02 lu0 = -1.054235903e-08 wu0 = -7.224255757e-09 pu0 = 3.167014752e-14
+ ua = -7.120310571e-10 lua = -2.898179157e-16 wua = -1.762999766e-17 pua = 1.124282282e-21
+ ub = 1.681817490e-18 lub = -6.022976162e-25 wub = -6.294868754e-25 pub = 1.505099045e-30
+ uc = -1.009067134e-10 luc = 9.029216596e-16 wuc = 5.270041644e-16 puc = -2.851051906e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.132572898e+00 la0 = 1.239921970e-06 wa0 = 1.075925533e-06 pa0 = -4.953361070e-12
+ ags = 2.585609582e-01 lags = 8.551777222e-07 wags = 3.059199105e-07 pags = -1.801789919e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.102384766e-24 lb0 = 2.447535939e-29 wb0 = 2.985245131e-29 pb0 = -1.197317938e-34
+ b1 = 0.0
+ keta = -1.001039642e-02 lketa = 2.450063773e-08 wketa = -1.829058468e-09 pketa = 4.463077187e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.589338897e-01 lpclm = 3.414210306e-06 wpclm = 1.042626713e-07 ppclm = -4.584614645e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 5.644443467e-03 lpdiblc2 = -1.116330436e-08 wpdiblc2 = -1.218471611e-08 ppdiblc2 = 5.617856901e-14
+ pdiblcb = 7.175821553e+00 lpdiblcb = -2.888095427e-05 wpdiblcb = -3.522592938e-05 ppdiblcb = 1.412836644e-10
+ drout = 0.56
+ pscbe1 = 3.047520763e+08 lpscbe1 = 1.975849033e+03 wpscbe1 = 1.394668907e+03 ppscbe1 = -5.563398338e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.570787832e-01 lkt1 = 1.684211460e-07 wkt1 = 1.242511916e-07 pkt1 = -5.386311418e-13
+ kt2 = -6.229710310e-02 lkt2 = 8.296108759e-08 wkt2 = 6.460144762e-08 pkt2 = -2.654721991e-13
+ at = 140000.0
+ ute = -2.359564205e+00 lute = 2.730163829e-06 wute = 1.567110738e-06 pute = -7.261293241e-12
+ ua1 = -4.790871812e-10 lua1 = 5.082008527e-15 wua1 = 2.470671323e-15 pua1 = -1.572461744e-20
+ ub1 = -1.856647873e-19 lub1 = -3.342840767e-24 wub1 = -9.084075536e-25 pub1 = 1.139602532e-29
+ uc1 = 2.750969333e-11 luc1 = -6.243490604e-17 wuc1 = -7.044317699e-17 puc1 = 4.589315736e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.21 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.849407657e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.954374892e-08 wvth0 = 1.493480423e-07 pvth0 = -3.085565420e-13
+ k1 = 5.392674576e-01 lk1 = 1.850575561e-08 wk1 = 2.170952134e-09 pk1 = 1.158792742e-13
+ k2 = -1.852913375e-02 lk2 = -2.963066067e-08 wk2 = -3.402362434e-08 pk2 = 2.932661985e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.297747128e+00 ldsub = -2.958945854e-06 wdsub = -2.133514529e-06 pdsub = 8.557070202e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.066412011e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.037156588e-08 wvoff = 4.090666117e-10 pvoff = -2.649953500e-14
+ nfactor = 3.954593718e+00 lnfactor = -2.419128404e-06 wnfactor = -6.202499164e-06 pnfactor = 1.256605759e-11
+ eta0 = 2.755029890e-01 leta0 = -7.841206513e-07 weta0 = -5.653813501e-07 peta0 = 2.267623603e-12
+ etab = -2.409114178e-01 letab = 6.854891218e-07 wetab = 4.942641983e-07 petab = -1.982387927e-12
+ u0 = 3.154354951e-02 lu0 = -2.694912393e-09 wu0 = 5.497287590e-09 pu0 = -1.935324044e-14
+ ua = -7.382552809e-10 lua = -1.846381661e-16 wua = 4.229457105e-16 pua = -6.427726000e-22
+ ub = 1.498593399e-18 lub = 1.325750035e-25 wub = 8.635602547e-26 pub = -1.365993640e-30
+ uc = 1.656480202e-10 luc = -1.661723340e-16 wuc = -3.137303798e-16 puc = 5.209544339e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.129692282e+00 la0 = -2.759310497e-06 wa0 = -2.673971892e-06 pa0 = 1.008667502e-11
+ ags = 4.749010050e-01 lags = -1.251590900e-08 wags = -7.389281037e-07 pags = 2.388871869e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.063517077e-24 lb0 = -1.228711140e-29 wb0 = -1.498651722e-29 pb0 = 6.010771345e-35
+ b1 = 0.0
+ keta = -1.066710308e-02 lketa = 2.713454760e-08 wketa = 2.573665998e-08 pketa = -6.592942575e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.025958054e-01 lpclm = -4.422795344e-07 wpclm = -3.731686384e-07 ppclm = 1.456413348e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 3.040775976e-04 lpdiblc2 = 1.025576030e-08 wpdiblc2 = 5.269413998e-09 ppdiblc2 = -1.382621168e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.826353960e+08 lpscbe1 = 5.916130450e+01 wpscbe1 = 7.446205589e+01 ppscbe1 = -2.683311812e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.952770924e-01 lkt1 = -7.945221035e-08 wkt1 = -5.698178526e-08 pkt1 = 1.882555444e-13
+ kt2 = -4.019920264e-02 lkt2 = -5.668862200e-09 wkt2 = -7.267174950e-09 pkt2 = 2.277746618e-14
+ at = 1.624029876e+05 lat = -8.985358906e-02 wat = 7.609535152e-03 pat = -3.052021705e-8
+ ute = -1.524983364e+00 lute = -6.171613213e-07 wute = -1.204123426e-06 pute = 3.853533948e-12
+ ua1 = 1.240370863e-09 lua1 = -1.814369724e-15 wua1 = -3.515337799e-15 pua1 = 8.283984142e-21
+ ub1 = -1.494323346e-18 lub1 = 1.905908658e-24 wub1 = 3.472993146e-24 pub1 = -6.176835269e-30
+ uc1 = 3.099794454e-12 luc1 = 3.546797465e-17 wuc1 = 1.804397813e-17 puc1 = 1.040285306e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.22 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.395544222e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.027262686e-08 wvth0 = -1.494186265e-07 pvth0 = 2.921992927e-13
+ k1 = 4.308356169e-01 lk1 = 2.365389830e-07 wk1 = 5.829737078e-07 pk1 = -1.051990776e-12
+ k2 = 3.908106057e-03 lk2 = -7.474714835e-08 wk2 = -1.794111518e-07 pk2 = 3.216698247e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.504620890e+00 ldsub = 2.676016523e-06 wdsub = 6.847680532e-06 pdsub = -9.502191090e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.444723420e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.425575203e-08 wvoff = 4.836491656e-08 pvoff = -1.229284867e-13
+ nfactor = 2.483487148e+00 lnfactor = 5.389520924e-07 wnfactor = 1.945379431e-06 pnfactor = -3.817582616e-12
+ eta0 = -2.276647030e-01 leta0 = 2.276418994e-07 weta0 = 1.116196192e-06 peta0 = -1.113668975e-12
+ etab = 7.880261914e-02 letab = 4.261261229e-08 wetab = -3.883071430e-07 petab = -2.077258298e-13
+ u0 = 3.294036187e-02 lu0 = -5.503603136e-09 wu0 = -1.632691007e-11 pu0 = -8.266541594e-15
+ ua = -3.258335162e-10 lua = -1.013930077e-15 wua = 6.515721262e-16 pua = -1.102491396e-21
+ ub = 9.565581684e-19 lub = 1.222491857e-24 wub = -1.030081871e-24 pub = 8.789240515e-31
+ uc = 1.513538305e-10 luc = -1.374297776e-16 wuc = -2.837677361e-16 puc = 4.607059694e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.398416014e+04 lvsat = 3.220442657e-02 wvsat = 5.922231393e-02 pvsat = -1.190833997e-7
+ a0 = -5.297877537e-01 la0 = 2.588334725e-06 wa0 = 7.872824655e-06 pa0 = -1.112067582e-11
+ ags = -2.734445773e-01 lags = 1.492246911e-06 wags = 7.758566726e-07 pags = -6.570361526e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.127034153e-24 lb0 = 6.193120344e-30 wb0 = 2.997303444e-29 pb0 = -3.029632359e-35
+ b1 = 0.0
+ keta = 9.607402992e-02 lketa = -1.874990283e-07 wketa = -1.255764835e-07 pketa = 2.383289247e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.242457111e+00 lpclm = -1.728903690e-06 wpclm = -3.261264820e-06 ppclm = 7.263756717e-12
+ pdiblc1 = 2.176329998e-01 lpdiblc1 = 3.465931508e-07 wpdiblc1 = -1.755111152e-07 ppdiblc1 = 3.529152932e-13
+ pdiblc2 = 3.176976609e-03 lpdiblc2 = 4.478975193e-09 wpdiblc2 = 9.421220314e-09 ppdiblc2 = -2.217460570e-14
+ pdiblcb = -5.031030115e-02 lpdiblcb = 5.089359921e-08 wpdiblcb = 6.778458428e-10 ppdiblcb = -1.363002931e-15
+ drout = 8.632358000e-01 ldrout = -6.097423013e-07 wdrout = -8.881784197e-22
+ pscbe1 = 5.779093808e+08 lpscbe1 = 4.708215096e+02 wpscbe1 = 1.705428261e+03 ppscbe1 = -3.547855193e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.347553610e-06 lalpha0 = 1.885625351e-11 walpha0 = 2.703506138e-11 palpha0 = -5.436172294e-17
+ alpha1 = 1.088945405e+00 lalpha1 = -4.804680759e-07 walpha1 = -1.337024352e-06 palpha1 = 2.688469848e-12
+ beta0 = 7.299595476e+00 lbeta0 = 1.319156957e-05 wbeta0 = 1.701667357e-05 pbeta0 = -3.421688898e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.694232834e-01 lkt1 = 6.963991258e-08 wkt1 = -5.954838544e-08 pkt1 = 1.934164281e-13
+ kt2 = -7.353752963e-02 lkt2 = 6.136737898e-08 wkt2 = 7.541524850e-08 pkt2 = -1.434791934e-13
+ at = 1.790757332e+05 lat = -1.233789125e-01 wat = -4.040650703e-02 pat = 6.602976834e-8
+ ute = -3.309734439e+00 lute = 2.971591154e-06 wute = 3.781460001e-06 pute = -6.171407408e-12
+ ua1 = -2.606269164e-09 lua1 = 5.920400189e-15 wua1 = 5.941249108e-15 pua1 = -1.073118842e-20
+ ub1 = 5.839796610e-19 lub1 = -2.273113932e-24 wub1 = 1.758326663e-25 pub1 = 4.530488623e-31
+ uc1 = -1.056356365e-10 luc1 = 2.541116569e-16 wuc1 = 6.108105077e-16 puc1 = -1.087898108e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.23 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.543335376e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.586745012e-08 wvth0 = 3.396081825e-07 pvth0 = -2.021021594e-13
+ k1 = 1.003286618e+00 lk1 = -3.420864745e-07 wk1 = -1.645208167e-06 pk1 = 1.200224268e-12
+ k2 = -1.865169406e-01 lk2 = 1.177318229e-07 wk2 = 5.358420685e-07 pk2 = -4.012981169e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.906612386e+00 ldsub = -7.720103144e-07 wdsub = -4.968312856e-06 pdsub = 2.441249603e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-7.604303952e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.275059435e-08 wvoff = -1.502504314e-07 pvoff = 7.782912636e-14
+ nfactor = 3.414547571e+00 lnfactor = -4.021507483e-07 wnfactor = -4.348498945e-06 pnfactor = 2.544181532e-12
+ eta0 = -5.055270701e-01 leta0 = 5.085012900e-07 weta0 = 2.913301718e-08 peta0 = -1.488073731e-14
+ etab = 2.443880222e-01 letab = -1.247587949e-07 wetab = -1.198184333e-06 petab = 6.108866954e-13
+ u0 = 2.733751508e-02 lu0 = 1.596759531e-10 wu0 = -2.386776792e-09 pu0 = -5.870524040e-15
+ ua = -1.156606155e-09 lua = -1.741967238e-16 wua = -5.961733011e-16 pua = 1.587122137e-22
+ ub = 2.013280681e-18 lub = 1.543715351e-25 wub = 3.115756508e-25 pub = -4.772045880e-31
+ uc = -6.064487983e-11 luc = 7.685555085e-17 wuc = 3.891609163e-16 puc = -2.194808914e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.514605742e+04 lvsat = 2.092213707e-02 wvsat = -1.906577960e-01 pvsat = 1.334919171e-7
+ a0 = 2.573307362e+00 la0 = -5.482303741e-07 wa0 = -6.325869750e-06 pa0 = 3.231165706e-12
+ ags = 1.057839332e+00 lags = 1.466037740e-07 wags = 7.284138074e-07 pags = -6.090815686e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.784463315e-01 lketa = 8.998230979e-08 wketa = 3.211334837e-07 pketa = -2.131992561e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.414364367e+00 lpclm = 9.565742645e-07 wpclm = 8.107120189e-06 ppclm = -4.227247693e-12
+ pdiblc1 = -3.233753597e-01 lpdiblc1 = 8.934368265e-07 wpdiblc1 = 3.086027705e-06 ppdiblc1 = -2.943802485e-12
+ pdiblc2 = 9.495128030e-03 lpdiblc2 = -1.907323810e-09 wpdiblc2 = -1.151446740e-08 ppdiblc2 = -1.013105651e-15
+ pdiblcb = 2.562060230e-02 lpdiblcb = -2.585629497e-08 wpdiblcb = -1.355691686e-09 ppdiblcb = 6.924683333e-16
+ drout = -2.892491878e-01 ldrout = 5.551733895e-07 wdrout = -5.978030981e-07 pdrout = 6.042510023e-13
+ pscbe1 = 1.292670842e+09 lpscbe1 = -2.516493687e+02 wpscbe1 = -3.648064366e+03 ppscbe1 = 1.863380205e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.352678562e-05 lalpha0 = -1.437266833e-11 walpha0 = -7.726609104e-11 palpha0 = 5.106442172e-17
+ alpha1 = 3.721091892e-01 lalpha1 = 2.440999357e-07 walpha1 = 2.674048704e-06 palpha1 = -1.365866641e-12
+ beta0 = 3.312283359e+01 lbeta0 = -1.291019799e-05 wbeta0 = -6.407971352e-05 pbeta0 = 4.775420374e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.240128802e-01 lkt1 = 2.373971274e-08 wkt1 = 2.713191202e-07 pkt1 = -1.410198144e-13
+ kt2 = 1.032328220e-02 lkt2 = -2.339795556e-08 wkt2 = -1.302520870e-07 pkt2 = 6.440647002e-14
+ at = 4.954612963e+04 lat = 7.547797404e-03 wat = 1.027532631e-01 pat = -7.867412304e-8
+ ute = 1.078885978e+00 lute = -1.464364923e-06 wute = -6.278721734e-06 pute = 3.997283446e-12
+ ua1 = 5.529613698e-09 lua1 = -2.303236305e-15 wua1 = -9.514522320e-15 pua1 = 4.891288959e-21
+ ub1 = -1.380475416e-18 lub1 = -2.874702419e-25 wub1 = -2.768687004e-24 pub1 = 3.429328122e-30
+ uc1 = 4.034149045e-10 luc1 = -2.604295032e-16 wuc1 = -1.409192782e-15 puc1 = 9.538929368e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.24 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.680040254e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.327244365e-08 wvth0 = -1.342643521e-07 pvth0 = 3.994529703e-14
+ k1 = -9.599558968e-02 lk1 = 2.194114872e-07 wk1 = 1.338287641e-06 pk1 = -3.237036211e-13
+ k2 = 1.855877311e-01 lk2 = -7.233403394e-08 wk2 = -4.859201458e-07 pk2 = 1.206037176e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.000602814e-01 ldsub = 4.859400894e-08 wdsub = -6.486766524e-07 pdsub = 2.348399052e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.399062768e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.301468342e-10 wvoff = 1.834511416e-08 pvoff = -8.287117955e-15
+ nfactor = 2.100585880e+00 lnfactor = 2.690024878e-07 wnfactor = 1.253257892e-06 pnfactor = -3.171174356e-13
+ eta0 = 0.49
+ etab = 2.143669139e-03 letab = -1.023770813e-09 wetab = -8.006802879e-09 petab = 2.960675575e-15
+ u0 = 3.841614930e-02 lu0 = -5.499135301e-09 wu0 = -2.132978318e-08 pu0 = 3.805298420e-15
+ ua = -8.244069547e-10 lua = -3.438794247e-16 wua = -7.543233911e-16 pua = 2.394930655e-22
+ ub = 2.052005131e-18 lub = 1.345916279e-25 wub = -3.208321031e-25 pub = -1.541795610e-31
+ uc = 1.741587971e-10 luc = -4.307888005e-17 wuc = -2.802302278e-16 puc = 1.224347335e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.042416423e+05 lvsat = 6.060519664e-03 wvsat = -4.539936912e-02 pvsat = 5.929594623e-8
+ a0 = 1.5
+ ags = 2.727358896e+00 lags = -7.061634462e-07 wags = -9.480701297e-07 pags = 2.472429557e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.763841729e-02 lketa = -1.017503471e-08 wketa = -1.407424350e-07 pketa = 2.272049684e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.358960122e-01 lpclm = 6.256576657e-08 wpclm = 4.227082817e-07 ppclm = -3.021576722e-13
+ pdiblc1 = 1.872845312e+00 lpdiblc1 = -2.283619457e-07 wpdiblc1 = -2.930628606e-06 ppdiblc1 = 1.294213259e-13
+ pdiblc2 = 9.203791952e-03 lpdiblc2 = -1.758513420e-09 wpdiblc2 = -2.794247220e-08 ppdiblc2 = 7.378089205e-15
+ pdiblcb = -3.266701514e-01 lpdiblcb = 1.540888900e-07 wpdiblcb = 1.475749867e-06 ppdiblcb = -7.537923717e-13
+ drout = 5.865718156e-01 ldrout = 1.078162825e-07 wdrout = 1.195606196e-06 pdrout = -3.117973575e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.592623138e-05 lalpha0 = 5.779380403e-12 walpha0 = 5.524643575e-11 palpha0 = -1.662112180e-17
+ alpha1 = 0.85
+ beta0 = -4.625052572e+00 lbeta0 = 6.370893794e-06 wbeta0 = 6.213664633e-05 pbeta0 = -1.671534584e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.405920253e-01 lkt1 = -1.887049208e-08 wkt1 = -2.107395881e-07 pkt1 = 1.052090250e-13
+ kt2 = -3.085713183e-02 lkt2 = -2.363576601e-09 wkt2 = -7.730641724e-08 pkt2 = 3.736256315e-14
+ at = 9.628588818e+04 lat = -1.632621690e-02 wat = -7.160444954e-02 pat = 1.038535556e-8
+ ute = -2.438414063e+00 lute = 3.322226955e-07 wute = 4.942141822e-07 pute = 5.377626013e-13
+ ua1 = 1.384509975e-09 lua1 = -1.859753549e-16 wua1 = -5.053915635e-15 pua1 = 2.612873513e-21
+ ub1 = -3.941920592e-18 lub1 = 1.020880094e-24 wub1 = 1.233486838e-23 pub1 = -4.285356519e-30
+ uc1 = -3.437286223e-10 luc1 = 1.212009503e-16 wuc1 = 1.148336553e-15 puc1 = -3.524572421e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.25 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {7.730160506e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.065810965e-08 wvth0 = -5.209818835e-07 pvth0 = 1.407958152e-13
+ k1 = 4.371245774e-01 lk1 = 8.038121129e-08 wk1 = -2.185173437e-08 pk1 = 3.100168605e-14
+ k2 = 5.507251898e-04 lk2 = -2.407897333e-08 wk2 = 1.231549536e-07 pk2 = -3.823454132e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 9.846145802e-01 ldsub = -1.299281684e-07 wdsub = -2.837501014e-07 pdsub = 1.396721697e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = -7.794471313e-03 lcdscd = 3.440933396e-09 wcdscd = 6.454645644e-08 pcdscd = -1.683281219e-14
+ cit = 0.0
+ voff = {-2.649240481e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.247273768e-08 wvoff = 6.382217716e-07 pvoff = -1.699422719e-13
+ nfactor = -9.830844703e-01 lnfactor = 1.073180544e-06 wnfactor = 1.681925887e-05 pnfactor = -4.376512567e-12
+ eta0 = 1.577656670e+00 leta0 = -2.836456324e-07 weta0 = 7.112806273e-07 peta0 = -1.854920297e-13
+ etab = -4.029506008e-02 letab = 1.004365563e-08 wetab = 5.130479682e-07 petab = -1.329231140e-13
+ u0 = -2.933691754e-02 lu0 = 1.216991599e-08 wu0 = 1.826920525e-08 pu0 = -6.521563375e-15
+ ua = -7.727338474e-09 lua = 1.456308474e-15 wua = 9.228952702e-15 pua = -2.364005574e-21
+ ub = 7.940176805e-18 lub = -1.400961110e-24 wub = -1.411045937e-23 pub = 3.441962174e-30
+ uc = -2.734310462e-10 luc = 7.364628480e-17 wuc = 1.121591051e-15 puc = -2.431406306e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.483384794e+05 lvsat = -5.439318103e-03 wvsat = 1.568731938e-01 pvsat = 6.546093629e-9
+ a0 = 1.5
+ ags = -3.334127560e+00 lags = 8.745873606e-07 wags = -6.588169051e-12 pags = 1.256930421e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.387875616e-02 lketa = -9.194567721e-09 wketa = -7.030020982e-08 pketa = 4.350150714e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.294973822e-01 lpclm = 1.207723970e-08 wpclm = -8.179378332e-08 ppclm = -1.705905967e-13
+ pdiblc1 = 2.619177152e+00 lpdiblc1 = -4.229948409e-07 wpdiblc1 = -8.713837152e-06 ppdiblc1 = 1.637601150e-12
+ pdiblc2 = -1.965367562e-02 lpdiblc2 = 5.767110119e-09 wpdiblc2 = 1.839232551e-08 ppdiblc2 = -4.705377350e-15
+ pdiblcb = 1.285093666e+00 lpdiblcb = -2.662365489e-07 wpdiblcb = -5.326361177e-06 ppdiblcb = 1.020102959e-12
+ drout = 3.561772454e-01 ldrout = 1.678999609e-07 wdrout = 5.776671875e-06 pdrout = -1.506475152e-12
+ pscbe1 = 7.823053059e+08 lpscbe1 = 4.614528506e+00 wpscbe1 = 1.188003750e+02 ppscbe1 = -3.098147460e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.184899916e-05 lalpha0 = -1.464010867e-12 walpha0 = 1.051022245e-12 palpha0 = -2.487716688e-18
+ alpha1 = 2.040839624e+00 lalpha1 = -3.105543021e-07 walpha1 = -3.443827214e-06 palpha1 = 8.981019240e-13
+ beta0 = 7.330784214e+00 lbeta0 = 3.252978942e-06 wbeta0 = 7.255437756e-05 pbeta0 = -1.943214430e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.361396470e-01 lkt1 = 6.046990006e-09 wkt1 = 2.963136104e-07 pkt1 = -2.702335043e-14
+ kt2 = -2.296425315e-02 lkt2 = -4.421928863e-09 wkt2 = 1.096797691e-07 pkt2 = -1.140081644e-14
+ at = 1.298124945e+05 lat = -2.506948646e-02 wat = -7.277514404e-01 pat = 1.814993047e-7
+ ute = 2.688182574e+00 lute = -1.004721935e-06 wute = -3.999067216e-07 pute = 7.709368153e-13
+ ua1 = 6.015080865e-09 lua1 = -1.393563415e-15 wua1 = 8.524450261e-15 pua1 = -9.281742155e-22
+ ub1 = -2.525137353e-18 lub1 = 6.514028599e-25 wub1 = -1.383568890e-23 pub1 = 2.539558431e-30
+ uc1 = 3.711290816e-10 luc1 = -6.522393088e-17 wuc1 = -1.686458139e-15 puc1 = 3.868175264e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.26 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.149419683e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.142118778e-08 wvth0 = 4.538638783e-07 pvth0 = -4.519110833e-14
+ k1 = 6.685934923e-01 lk1 = 3.622018288e-08 wk1 = 6.896679366e-07 pk1 = -1.047463059e-13
+ k2 = -9.081029267e-02 lk2 = -6.648570177e-09 wk2 = -9.400709982e-08 pk2 = 3.196938201e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.380909432e-01 ldsub = -6.580509818e-09 wdsub = 3.486673228e-07 pdsub = 1.901577900e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 3.572544955e-02 lcdscd = -4.862058226e-09 wcdscd = -9.738132631e-08 pcdscd = 1.406074177e-14
+ cit = 0.0
+ voff = {1.451800107e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.576937528e-08 wvoff = -9.462980199e-07 pvoff = 1.323619210e-13
+ nfactor = 1.284791319e+01 lnfactor = -1.565580175e-06 wnfactor = -3.858105295e-05 pnfactor = 6.193091324e-12
+ eta0 = 5.743312101e-01 leta0 = -9.222518117e-08 weta0 = -1.658919380e-06 peta0 = 2.667089490e-13
+ etab = 1.845252169e-01 letab = -3.284890573e-08 wetab = -6.815885125e-07 petab = 9.499680166e-14
+ u0 = 2.268845522e-01 lu0 = -3.671355334e-08 wu0 = -5.877601969e-07 pu0 = 1.091003621e-13
+ ua = 2.167070205e-08 lua = -4.152426084e-15 wua = -6.610658633e-14 pua = 1.200896058e-20
+ ub = -1.779112800e-17 lub = 3.508211608e-24 wub = 5.681220109e-23 pub = -1.008908852e-29
+ uc = 6.326668275e-10 luc = -9.922450413e-17 wuc = -1.656868318e-15 puc = 2.869505187e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.186456878e+05 lvsat = 6.457612321e-02 wvsat = 9.439076799e-01 pvsat = -1.436090678e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.981917596e-01 lketa = -1.397519084e-07 wketa = -3.237749247e-06 pketa = 6.086550827e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.125584191e+00 lpclm = -4.832197783e-07 wpclm = -6.816511825e-06 ppclm = 1.114299320e-12
+ pdiblc1 = 8.154212105e-01 lpdiblc1 = -7.886345980e-08 wpdiblc1 = -1.325803508e-06 ppdiblc1 = 2.280677630e-13
+ pdiblc2 = 1.563707289e-02 lpdiblc2 = -9.658706263e-10 wpdiblc2 = -2.091144689e-08 ppdiblc2 = 2.793232172e-15
+ pdiblcb = -1.032864742e+00 lpdiblcb = 1.759974640e-07 wpdiblcb = 2.688250257e-06 ppdiblcb = -5.089726980e-13
+ drout = 5.500528586e+00 ldrout = -8.135702539e-07 wdrout = -1.445156816e-05 pdrout = 2.352789852e-12
+ pscbe1 = 8.766256060e+08 lpscbe1 = -1.338046427e+01 wpscbe1 = -2.464091656e+02 ppscbe1 = 3.869539281e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.639295687e-05 lalpha0 = -4.238794384e-12 walpha0 = -7.623987860e-11 palpha0 = 1.225830512e-17
+ alpha1 = -1.928625788e+00 lalpha1 = 4.467641260e-07 walpha1 = 8.035596834e-06 palpha1 = -1.292011473e-12
+ beta0 = 8.076986596e+01 lbeta0 = -1.075816971e-05 wbeta0 = -1.863261607e-04 pbeta0 = 2.995863807e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.289936741e-01 lkt1 = 8.099803842e-08 wkt1 = 1.382438739e-06 pkt1 = -2.342408193e-13
+ kt2 = -1.346858683e-01 lkt2 = 1.689299121e-08 wkt2 = 3.059864447e-07 pkt2 = -4.885338186e-14
+ at = -3.104658499e+05 lat = 5.892945775e-02 wat = 1.349315715e+00 pat = -2.147760296e-7
+ ute = -2.661733750e+01 lute = 4.586361017e-06 wute = 7.316094682e-05 pute = -1.326344419e-11
+ ua1 = -3.216063602e-08 lua1 = 5.889828907e-15 wua1 = 9.293740757e-14 pua1 = -1.703298469e-20
+ ub1 = 1.915179126e-17 lub1 = -3.484251643e-24 wub1 = -5.333890397e-23 pub1 = 1.007621882e-29
+ uc1 = -5.103039945e-10 luc1 = 1.029411600e-16 wuc1 = 1.901417078e-15 puc1 = -2.976988347e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.27 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.037705701e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.743443722e-07 wvth0 = 3.099505687e-08 pvth0 = -6.202354501e-13
+ k1 = 5.345769059e-01 lk1 = 3.379922632e-07 wk1 = 1.051759441e-08 pk1 = -2.104653309e-13
+ k2 = -2.169276183e-02 lk2 = -1.972361156e-07 wk2 = -1.100274930e-08 pk2 = 2.201736616e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.079585345e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.422912971e-08 wvoff = 8.126087911e-09 pvoff = -1.626094062e-13
+ nfactor = 3.264920145e+00 lnfactor = -1.648829025e-05 wnfactor = -1.502249661e-06 pnfactor = 3.006119649e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.143810506e-02 lu0 = -7.704253888e-09 wu0 = 3.652512495e-10 pu0 = -7.308964590e-15
+ ua = -8.534025596e-10 lua = 2.954131897e-15 wua = 2.382679590e-16 pua = -4.767929139e-21
+ ub = 1.727672372e-18 lub = -5.477800018e-24 wub = -3.702443845e-25 pub = 7.408881147e-30
+ uc = 4.962252348e-11 luc = 4.272198059e-16 wuc = -1.681934124e-17 puc = 3.365682383e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.323342844e+00 la0 = 2.446141610e-06 wa0 = 7.826910202e-08 pa0 = -1.566226251e-12
+ ags = 3.723302380e-01 lags = 4.200816687e-07 wags = 1.263331569e-08 pags = -2.528025767e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.271091167e-25 lb0 = 5.271659707e-29
+ b1 = 7.618685315e-24 lb1 = -1.524558814e-28 wb1 = -1.441403454e-29 pb1 = 2.884361607e-34
+ keta = -1.574673177e-02 lketa = 2.018854536e-07 wketa = 1.783608855e-08 pketa = -3.569141510e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.075926543e-01 lpclm = 3.824534545e-06 wpclm = 3.458669416e-07 ppclm = -6.921069353e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.941906546e-03 lpdiblc2 = -9.592555392e-09 wpdiblc2 = 8.223638722e-10 ppdiblc2 = -1.645614746e-14
+ pdiblcb = 5.969894081e-01 lpdiblcb = -6.220564959e-05 wpdiblcb = 1.942890293e-22 ppdiblcb = 9.769962617e-27
+ drout = 0.56
+ pscbe1 = 8.872089763e+08 lpscbe1 = -1.874874501e+03 wpscbe1 = -4.113786519e+02 ppscbe1 = 8.232010169e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.853100699e-01 lkt1 = -6.209332904e-07 wkt1 = -7.776978851e-08 pkt1 = 1.556234595e-12
+ kt2 = -4.591286303e-02 lkt2 = 9.707634562e-08 wkt2 = -1.341757989e-09 pkt2 = 2.684963198e-14
+ at = 140000.0
+ ute = -1.652906658e+00 lute = -2.749348768e-06 wute = -4.808457460e-07 pute = 9.622101323e-12
+ ua1 = 6.638467717e-10 lua1 = -6.662926814e-15 wua1 = -7.997223987e-16 pua1 = 1.600307378e-20
+ ub1 = -1.028574077e-18 lub1 = 1.207478996e-23 wub1 = 9.696941880e-25 pub1 = -1.940434288e-29
+ uc1 = 1.316378282e-11 luc1 = 4.009259381e-17 wuc1 = 8.188837255e-18 puc1 = -1.638650699e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.28 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.5224777+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55146741
+ k2 = -0.031549252
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.44095
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0310531
+ ua = -7.0577558e-10
+ ub = 1.45393e-18
+ uc = 7.0972e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.445584
+ ags = 0.393323
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.1073e-24
+ b1 = 0.0
+ keta = -0.0056579
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0024625373
+ pdiblcb = -2.5116166
+ drout = 0.56
+ pscbe1 = 793515780.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31634
+ kt2 = -0.041061662
+ at = 140000.0
+ ute = -1.7903
+ ua1 = 3.3088e-10
+ ub1 = -4.2516e-19
+ uc1 = 1.5167332e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.29 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.101215713e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.898230280e-8
+ k1 = 5.483036418e-01 lk1 = 2.534426967e-8
+ k2 = -2.793528414e-02 lk2 = -2.895072312e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.077968391e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.641064876e-8
+ nfactor = 2.592246875e+00 lnfactor = -1.212006887e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.100206275e-02 lu0 = 4.088485026e-10
+ ua = -7.181273269e-10 lua = 9.894720127e-17
+ ub = 1.464147477e-18 lub = -8.185002439e-26
+ uc = 8.132584406e-11 luc = -8.294242903e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.504616754e+00 la0 = -4.728987572e-7
+ ags = 3.643448806e-01 lags = 2.321375129e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.220282334e-24 lb0 = -1.692664930e-29
+ b1 = 0.0
+ keta = -1.064286581e-02 lketa = 3.993349433e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.228809427e-01 lpclm = 3.255679101e-06 wpclm = -1.110223025e-22 ppclm = 1.332267630e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.431095396e-03 lpdiblc2 = 8.262660361e-9
+ pdiblcb = -5.004938362e+00 lpdiblcb = 1.997346706e-05 ppdiblcb = 1.421085472e-26
+ drout = 0.56
+ pscbe1 = 7.870140753e+08 lpscbe1 = 5.208376498e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.141140138e-01 lkt1 = -1.783189933e-8
+ kt2 = -3.995859458e-02 lkt2 = -8.836437064e-9
+ at = 140000.0
+ ute = -1.817673614e+00 lute = 2.192841674e-7
+ ua1 = 3.752452592e-10 lua1 = -3.554005973e-16
+ ub1 = -4.997826689e-19 lub1 = 5.977862313e-25
+ uc1 = 3.151175570e-12 luc1 = 9.625885770e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.30 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.365837650e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.151893317e-9
+ k1 = 5.400181503e-01 lk1 = 5.857560310e-8
+ k2 = -3.029414909e-02 lk2 = -1.948982062e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.064997501e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.120830236e-8
+ nfactor = 1.809834034e+00 lnfactor = 1.926083583e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.344445436e-02 lu0 = -9.387061600e-9
+ ua = -5.920050542e-10 lua = -4.069022443e-16
+ ub = 1.528454414e-18 lub = -3.397713864e-25
+ uc = 5.716331865e-11 luc = 1.396828961e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.205060620e+00 la0 = 7.285567913e-7
+ ags = 2.193873541e-01 lags = 8.135311311e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.118664669e-24 lb0 = 8.497510593e-30
+ b1 = 0.0
+ keta = -1.767633807e-03 lketa = 4.336838064e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.735579725e-01 lpclm = 6.133304993e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 2.126186139e-03 lpdiblc2 = 5.474800142e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.083836002e+08 lpscbe1 = -3.362482644e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.149808009e-01 lkt1 = -1.435540156e-8
+ kt2 = -4.271211613e-02 lkt2 = 2.207348643e-9
+ at = 1.650342857e+05 lat = -1.004071626e-1
+ ute = -1.941356718e+00 lute = 7.153506284e-7
+ ua1 = 2.480362285e-11 lua1 = 1.050145812e-15
+ ub1 = -2.933984465e-19 lub1 = -2.299767186e-25
+ uc1 = 9.339214374e-12 luc1 = 7.143995830e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.31 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.878870156e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.076684872e-8
+ k1 = 6.324218602e-01 lk1 = -1.272284831e-7
+ k2 = -5.813040379e-02 lk2 = 3.648293062e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.772314921e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.676314387e-8
+ nfactor = 3.156179117e+00 lnfactor = -7.811282609e-7
+ eta0 = 1.583043279e-01 leta0 = -1.574532464e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 3.293471619e-02 lu0 = -8.362087220e-9
+ ua = -1.005266535e-10 lua = -1.395160132e-15
+ ub = 6.003665738e-19 lub = 1.526414650e-24
+ uc = 5.322989950e-11 luc = 2.187755377e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.446262019e+04 lvsat = -8.973374201e-3
+ a0 = 2.192553109e+00 la0 = -1.257079281e-6
+ ags = -5.161411334e-03 lags = 1.265050645e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.237329338e-24 lb0 = -4.283033172e-30
+ b1 = 0.0
+ keta = 5.265098834e-02 lketa = -1.050873655e-07 wketa = 1.647987302e-23 pketa = -5.464378949e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.147456642e-01 lpclm = 7.828278159e-7
+ pdiblc1 = 1.569430821e-01 lpdiblc1 = 4.686275877e-7
+ pdiblc2 = 6.434736582e-03 lpdiblc2 = -3.188772769e-9
+ pdiblcb = -5.007590911e-02 lpdiblcb = 5.042228697e-8
+ drout = 8.632358000e-01 ldrout = -6.097423013e-7
+ pscbe1 = 1.167628731e+09 lpscbe1 = -7.559899069e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 8.893632000e-10 lalpha0 = 5.853526093e-14
+ alpha1 = 6.266162940e-01 lalpha1 = 4.491768287e-7
+ beta0 = 1.318378417e+01 lbeta0 = 1.359725332e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.900144956e-01 lkt1 = 1.365213013e-7
+ kt2 = -4.745972127e-02 lkt2 = 1.175376658e-8
+ at = 1.651035834e+05 lat = -1.005465055e-1
+ ute = -2.002144911e+00 lute = 8.375826746e-7
+ ua1 = -5.518470310e-10 lua1 = 2.209666873e-15
+ ub1 = 6.447807678e-19 lub1 = -2.116454348e-24
+ uc1 = 1.055762826e-10 luc1 = -1.220721912e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.32 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.717665141e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.982625921e-9
+ k1 = 4.343907494e-01 lk1 = 7.293859126e-8
+ k2 = -1.228327853e-03 lk2 = -2.103289110e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.886214874e-01 ldsub = 7.214840124e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.279980756e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.838092139e-9
+ nfactor = 1.910881874e+00 lnfactor = 4.776007576e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 6.938893904e-23 peta0 = 1.786765180e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.651219250e-02 lu0 = -1.870290187e-9
+ ua = -1.362756681e-09 lua = -1.193156915e-16
+ ub = 2.121020299e-18 lub = -1.064084691e-26
+ uc = 7.392291647e-11 luc = 9.613419190e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.218575020e+03 lvsat = 6.708225324e-2
+ a0 = 3.858874119e-01 la0 = 5.690731124e-7
+ ags = 1.309717248e+00 lags = -6.401029598e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.740171369e-02 lketa = 1.626022499e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.388993454e+00 lpclm = -5.051640103e-7
+ pdiblc1 = 7.437409158e-01 lpdiblc1 = -1.244994474e-07 wpdiblc1 = 8.881784197e-22
+ pdiblc2 = 5.513544990e-03 lpdiblc2 = -2.257645204e-9
+ pdiblcb = 2.515181822e-02 lpdiblcb = -2.561684662e-08 wpdiblcb = 1.214306433e-23 ppdiblcb = 2.168404345e-31
+ drout = -4.959632800e-01 ldrout = 7.641170999e-7
+ pscbe1 = 3.120813611e+07 lpscbe1 = 3.926881210e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.191024846e-06 lalpha0 = 3.284877457e-12 walpha0 = -1.482307658e-27 palpha0 = 7.411538288e-34
+ alpha1 = 1.296767412e+00 lalpha1 = -2.282025393e-7
+ beta0 = 1.096473529e+01 lbeta0 = 3.602708867e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.301935511e-01 lkt1 = -2.502347200e-8
+ kt2 = -3.471653443e-02 lkt2 = -1.126868269e-9
+ at = 8.507713903e+04 lat = -1.965689587e-2
+ ute = -1.092230678e+00 lute = -8.214589253e-8
+ ua1 = 2.239590862e-09 lua1 = -6.118794686e-16
+ ub1 = -2.337858579e-18 lub1 = 8.983557464e-25
+ uc1 = -8.386929930e-11 luc1 = 6.941675076e-17 wuc1 = 2.584939414e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.33 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.215768093e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.945977550e-8
+ k1 = 3.667703539e-01 lk1 = 1.074781426e-7
+ k2 = 1.756159980e-02 lk2 = -3.063052309e-08 pk2 = 1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 7.575464332e-02 ldsub = 1.297992051e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.335627272e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.995746010e-9
+ nfactor = 2.533949421e+00 lnfactor = 1.593465777e-7
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 3.104053217e-02 lu0 = -4.183302695e-9
+ ua = -1.085244136e-09 lua = -2.610652142e-16
+ ub = 1.941064728e-18 lub = 8.127793964e-26
+ uc = 7.725809959e-11 luc = -7.422229282e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.854301274e+04 lvsat = 2.656444100e-2
+ a0 = 1.5
+ ags = 2.399526108e+00 lags = -6.206694043e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.102885254e-02 lketa = -2.318523268e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.820641385e-01 lpclm = -4.191721304e-8
+ pdiblc1 = 8.594644286e-01 lpdiblc1 = -1.836093976e-7
+ pdiblc2 = -4.584242403e-04 lpdiblc2 = 7.927530709e-10 ppdiblc2 = 4.336808690e-31
+ pdiblcb = 1.836288000e-01 lpdiblcb = -1.065646702e-07 wpdiblcb = -1.110223025e-22
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.177411360e-06 lalpha0 = 3.196940107e-14
+ alpha1 = 0.85
+ beta0 = 1.686115330e+01 lbeta0 = 5.909010965e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.134635824e-01 lkt1 = 1.750969425e-8
+ kt2 = -5.758888667e-02 lkt2 = 1.055600904e-8
+ at = 7.152581445e+04 lat = -1.273506899e-2
+ ute = -2.267519941e+00 lute = 5.181754085e-7
+ ua1 = -3.630814747e-10 lua1 = 7.175291234e-16
+ ub1 = 3.233485706e-19 lub1 = -4.609516086e-25 pub1 = -1.925929944e-46
+ uc1 = 5.335421127e-11 luc1 = -6.750973096e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.34 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.826818720e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.316520387e-09 wvth0 = 2.945161824e-08 pvth0 = -7.680569715e-15
+ k1 = 4.295684749e-01 lk1 = 9.110127180e-8
+ k2 = 6.613024587e-03 lk2 = -2.777528795e-08 wk2 = 1.056231960e-07 pk2 = -2.754505078e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.864712740e-01 ldsub = -8.162434218e-08 wdsub = 7.366632614e-11 pdsub = -1.921114653e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 1.452502183e-02 lcdscd = -2.379677943e-09 wcdscd = -1.387778781e-23
+ cit = 0.0
+ voff = {-1.756724704e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.985885496e-09 wvoff = 3.801122780e-07 pvoff = -9.912796053e-14
+ nfactor = 2.349537676e+00 lnfactor = 2.074385790e-07 wnfactor = 7.181542241e-06 pnfactor = -1.872845675e-12
+ eta0 = 1.823610105e+00 leta0 = -3.477868449e-07 weta0 = 1.819289785e-14 peta0 = -4.744453275e-21
+ etab = 1.740475113e-01 letab = -4.555214553e-08 wetab = -1.068161729e-07 petab = 2.785616247e-14
+ u0 = -1.260304720e-02 lu0 = 7.198331796e-09 wu0 = -3.012400987e-08 pu0 = 7.855920038e-15
+ ua = -4.266324707e-09 lua = 5.685160635e-16 wua = -7.800637625e-16 pua = 2.034297084e-22
+ ub = 1.928304229e-18 lub = 8.460569905e-26 wub = 3.275467315e-24 pub = -8.541960192e-31
+ uc = 2.314608982e-10 luc = -4.095615398e-17 wuc = -3.385221194e-16 puc = 8.828182942e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.036146612e+05 lvsat = -2.952323392e-02 wvsat = -2.921749652e-01 pvsat = 7.619514047e-8
+ a0 = 1.5
+ ags = -3.334129838e+00 lags = 8.745877952e-07 wags = -5.551115123e-22 pags = -3.330669074e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.461768944e-01 lketa = -1.006885012e-07 wketa = -1.031283829e-06 pketa = 2.689443847e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.541814529e-02 lpclm = 9.042706182e-08 wpclm = 1.522984188e-06 ppclm = -3.971729544e-13
+ pdiblc1 = -3.939770822e-01 lpdiblc1 = 1.432706002e-7
+ pdiblc2 = -1.329380080e-02 lpdiblc2 = 4.140039583e-09 wpdiblc2 = 6.938893904e-24 ppdiblc2 = -1.734723476e-30
+ pdiblcb = -5.567066175e-01 lpdiblcb = 8.650444195e-8
+ drout = 2.353690284e+00 ldrout = -3.530234743e-7
+ pscbe1 = 8.233852396e+08 lpscbe1 = -6.098543103e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.221243171e-05 lalpha0 = -2.324237417e-12
+ alpha1 = 0.85
+ beta0 = 3.040830297e+01 lbeta0 = -2.942005877e-06 wbeta0 = 5.815762590e-06 pbeta0 = -1.516669463e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.821126062e-01 lkt1 = -1.674480144e-08 wkt1 = -1.491221177e-07 pkt1 = 3.888896058e-14
+ kt2 = 1.496186997e-02 lkt2 = -8.364212580e-9
+ at = -1.991836980e+05 lat = 5.786218192e-02 wat = 2.236831765e-01 pat = -5.833344087e-8
+ ute = 2.549898990e+00 lute = -7.381400046e-07 pute = 4.440892099e-28
+ ua1 = 8.962747083e-09 lua1 = -1.714516403e-15
+ ub1 = -7.309374636e-18 lub1 = 1.529555746e-24
+ uc1 = -2.120305980e-10 luc1 = 6.853354557e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.35 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {9.438398519e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.822040675e-08 wvth0 = -7.864796361e-07 pvth0 = 1.479876906e-13
+ k1 = 0.90707349
+ k2 = -5.494816598e-02 lk2 = -1.603027465e-08 wk2 = -1.977179316e-07 pk2 = 3.032818958e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587159132e-01 ldsub = -1.460792414e-11 wdsub = -1.718880943e-10 pdsub = 2.763719913e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-1.338146533e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -1.394644233e-7
+ nfactor = -5.293063660e+00 lnfactor = 1.665539917e-06 wnfactor = 1.388141850e-05 pnfactor = -3.151088267e-12
+ eta0 = 6.941612174e-04 leta0 = -3.607624990e-15 weta0 = -4.245009617e-14 peta0 = 6.825381162e-21
+ etab = -6.471290892e-02 wetab = 3.919119906e-8
+ u0 = 9.783655146e-03 lu0 = 2.927262402e-09 wu0 = 4.008083455e-08 pu0 = -5.538181410e-15
+ ua = -1.288698684e-09 lua = 4.267051525e-19 wua = 2.904393431e-16 pua = -8.072971326e-25
+ ub = 2.076034198e-18 lub = 5.642088919e-26 wub = -6.422810181e-25 pub = -1.067444857e-31
+ uc = 1.679025167e-11 wuc = 1.242048597e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.725145711e+04 lvsat = 4.314068933e-02 wvsat = 5.350051796e-01 pvsat = -8.161925064e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.253471759e+00 lketa = 2.045020667e-07 wketa = 2.406328935e-06 pketa = -3.869040041e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.932621135e+00 lpclm = -2.831394203e-07 wpclm = -3.366543787e-06 ppclm = 5.356805298e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 2.103262180e+01 lbeta0 = -1.153257169e-06 wbeta0 = -1.357011271e-05 pbeta0 = 2.181884142e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.698800600e-01 wkt1 = 5.471338693e-8
+ kt2 = -0.028878939
+ at = 3.365905563e+05 lat = -4.435604496e-02 wat = -5.219274119e-01 pat = 8.391862085e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.36 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.201533243e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.651258432e-8
+ k1 = 5.401360879e-01 lk1 = 2.267486609e-7
+ k2 = -2.750837745e-02 lk2 = -8.086107591e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.036634077e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.171973431e-8
+ nfactor = 2.470890729e+00 lnfactor = -5.991375219e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.163116234e-02 lu0 = -1.156748184e-8
+ ua = -7.274635940e-10 lua = 4.339942073e-16
+ ub = 1.531975917e-18 lub = -1.561760146e-24
+ uc = 4.073248872e-11 luc = 6.051163890e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.364712778e+00 la0 = 1.618296714e-6
+ ags = 3.790077061e-01 lags = 2.864602824e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.271091167e-25 lb0 = 5.271659707e-29
+ b1 = 0.0
+ keta = -6.319284829e-03 lketa = 1.323483028e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.521885355e-02 lpclm = 1.663325838e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.376575378e-03 lpdiblc2 = -1.829062036e-8
+ pdiblcb = 5.969894081e-01 lpdiblcb = -6.220564959e-05 wpdiblcb = -2.775557562e-22 ppdiblcb = -3.907985047e-26
+ drout = 0.56
+ pscbe1 = 6.697705843e+08 lpscbe1 = 2.476238630e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.264160867e-01 lkt1 = 2.016304145e-7
+ kt2 = -4.662206293e-02 lkt2 = 1.112679931e-7
+ at = 140000.0
+ ute = -1.907062593e+00 lute = 2.336511254e-6
+ ua1 = 2.411453223e-10 lua1 = 1.795661433e-15
+ ub1 = -5.160323004e-19 lub1 = 1.818426157e-24
+ uc1 = 1.749207647e-11 luc1 = -4.651996409e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.37 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.5224777+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55146741
+ k2 = -0.031549252
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.44095
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0310531
+ ua = -7.0577558e-10
+ ub = 1.45393e-18
+ uc = 7.0972e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.445584
+ ags = 0.393323
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.1073e-24
+ b1 = 0.0
+ keta = -0.0056579
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0024625373
+ pdiblcb = -2.5116166
+ drout = 0.56
+ pscbe1 = 793515780.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31634
+ kt2 = -0.041061662
+ at = 140000.0
+ ute = -1.7903
+ ua1 = 3.3088e-10
+ ub1 = -4.2516e-19
+ uc1 = 1.5167332e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.38 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.101215713e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.898230280e-8
+ k1 = 5.483036418e-01 lk1 = 2.534426967e-8
+ k2 = -2.793528414e-02 lk2 = -2.895072312e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.077968391e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.641064876e-8
+ nfactor = 2.592246875e+00 lnfactor = -1.212006887e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.100206275e-02 lu0 = 4.088485026e-10
+ ua = -7.181273269e-10 lua = 9.894720127e-17
+ ub = 1.464147477e-18 lub = -8.185002439e-26
+ uc = 8.132584406e-11 luc = -8.294242903e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.504616754e+00 la0 = -4.728987572e-7
+ ags = 3.643448806e-01 lags = 2.321375129e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.220282334e-24 lb0 = -1.692664930e-29
+ b1 = 0.0
+ keta = -1.064286581e-02 lketa = 3.993349433e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.228809427e-01 lpclm = 3.255679101e-06 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.431095396e-03 lpdiblc2 = 8.262660361e-9
+ pdiblcb = -5.004938362e+00 lpdiblcb = 1.997346706e-5
+ drout = 0.56
+ pscbe1 = 7.870140753e+08 lpscbe1 = 5.208376498e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.141140138e-01 lkt1 = -1.783189933e-8
+ kt2 = -3.995859458e-02 lkt2 = -8.836437064e-9
+ at = 140000.0
+ ute = -1.817673614e+00 lute = 2.192841674e-7
+ ua1 = 3.752452592e-10 lua1 = -3.554005973e-16
+ ub1 = -4.997826689e-19 lub1 = 5.977862313e-25
+ uc1 = 3.151175570e-12 luc1 = 9.625885770e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.39 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.365837650e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.151893317e-9
+ k1 = 5.400181503e-01 lk1 = 5.857560310e-8
+ k2 = -3.029414909e-02 lk2 = -1.948982062e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.064997501e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.120830236e-8
+ nfactor = 1.809834034e+00 lnfactor = 1.926083583e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.344445436e-02 lu0 = -9.387061600e-9
+ ua = -5.920050542e-10 lua = -4.069022443e-16
+ ub = 1.528454414e-18 lub = -3.397713864e-25
+ uc = 5.716331865e-11 luc = 1.396828961e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.205060620e+00 la0 = 7.285567913e-7
+ ags = 2.193873541e-01 lags = 8.135311311e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.118664669e-24 lb0 = 8.497510593e-30
+ b1 = 0.0
+ keta = -1.767633807e-03 lketa = 4.336838064e-09 wketa = -1.734723476e-24
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.735579725e-01 lpclm = 6.133304993e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 2.126186139e-03 lpdiblc2 = 5.474800142e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.083836002e+08 lpscbe1 = -3.362482644e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.149808009e-01 lkt1 = -1.435540156e-8
+ kt2 = -4.271211613e-02 lkt2 = 2.207348643e-9
+ at = 1.650342857e+05 lat = -1.004071626e-1
+ ute = -1.941356718e+00 lute = 7.153506284e-7
+ ua1 = 2.480362285e-11 lua1 = 1.050145812e-15
+ ub1 = -2.933984465e-19 lub1 = -2.299767186e-25
+ uc1 = 9.339214374e-12 luc1 = 7.143995830e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.40 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.878870156e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.076684872e-8
+ k1 = 6.324218602e-01 lk1 = -1.272284831e-7
+ k2 = -5.813040379e-02 lk2 = 3.648293062e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.772314921e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.676314387e-8
+ nfactor = 3.156179117e+00 lnfactor = -7.811282609e-7
+ eta0 = 1.583043279e-01 leta0 = -1.574532464e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 3.293471619e-02 lu0 = -8.362087220e-9
+ ua = -1.005266535e-10 lua = -1.395160132e-15
+ ub = 6.003665738e-19 lub = 1.526414650e-24
+ uc = 5.322989950e-11 luc = 2.187755377e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.446262019e+04 lvsat = -8.973374201e-3
+ a0 = 2.192553109e+00 la0 = -1.257079281e-6
+ ags = -5.161411334e-03 lags = 1.265050645e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.237329338e-24 lb0 = -4.283033172e-30
+ b1 = 0.0
+ keta = 5.265098834e-02 lketa = -1.050873655e-07 wketa = 2.428612866e-23 pketa = 4.336808690e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.147456642e-01 lpclm = 7.828278159e-7
+ pdiblc1 = 1.569430821e-01 lpdiblc1 = 4.686275877e-7
+ pdiblc2 = 6.434736582e-03 lpdiblc2 = -3.188772769e-9
+ pdiblcb = -5.007590911e-02 lpdiblcb = 5.042228697e-8
+ drout = 8.632358000e-01 ldrout = -6.097423013e-7
+ pscbe1 = 1.167628731e+09 lpscbe1 = -7.559899069e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 8.893632000e-10 lalpha0 = 5.853526093e-14
+ alpha1 = 6.266162940e-01 lalpha1 = 4.491768287e-7
+ beta0 = 1.318378417e+01 lbeta0 = 1.359725332e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.900144956e-01 lkt1 = 1.365213013e-7
+ kt2 = -4.745972127e-02 lkt2 = 1.175376658e-8
+ at = 1.651035834e+05 lat = -1.005465055e-1
+ ute = -2.002144911e+00 lute = 8.375826746e-7
+ ua1 = -5.518470310e-10 lua1 = 2.209666873e-15
+ ub1 = 6.447807678e-19 lub1 = -2.116454348e-24
+ uc1 = 1.055762826e-10 luc1 = -1.220721912e-16 wuc1 = -1.033975766e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.41 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.717665141e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.982625921e-9
+ k1 = 4.343907494e-01 lk1 = 7.293859126e-8
+ k2 = -1.228327853e-03 lk2 = -2.103289110e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.886214874e-01 ldsub = 7.214840124e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.279980756e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.838092139e-9
+ nfactor = 1.910881874e+00 lnfactor = 4.776007576e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -4.093947403e-22 peta0 = 7.285838599e-29
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.651219250e-02 lu0 = -1.870290187e-9
+ ua = -1.362756681e-09 lua = -1.193156915e-16
+ ub = 2.121020299e-18 lub = -1.064084691e-26
+ uc = 7.392291647e-11 luc = 9.613419190e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.218575020e+03 lvsat = 6.708225324e-2
+ a0 = 3.858874119e-01 la0 = 5.690731124e-7
+ ags = 1.309717248e+00 lags = -6.401029598e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.740171369e-02 lketa = 1.626022499e-08 wketa = -1.110223025e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.388993454e+00 lpclm = -5.051640103e-7
+ pdiblc1 = 7.437409158e-01 lpdiblc1 = -1.244994474e-7
+ pdiblc2 = 5.513544990e-03 lpdiblc2 = -2.257645204e-9
+ pdiblcb = 2.515181822e-02 lpdiblcb = -2.561684662e-08 wpdiblcb = -1.084202172e-23 ppdiblcb = 8.673617380e-30
+ drout = -4.959632800e-01 ldrout = 7.641170999e-7
+ pscbe1 = 3.120813611e+07 lpscbe1 = 3.926881210e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.191024846e-06 lalpha0 = 3.284877457e-12 walpha0 = 1.270549421e-27
+ alpha1 = 1.296767412e+00 lalpha1 = -2.282025393e-7
+ beta0 = 1.096473529e+01 lbeta0 = 3.602708867e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.301935511e-01 lkt1 = -2.502347200e-8
+ kt2 = -3.471653443e-02 lkt2 = -1.126868269e-9
+ at = 8.507713903e+04 lat = -1.965689587e-2
+ ute = -1.092230678e+00 lute = -8.214589253e-8
+ ua1 = 2.239590862e-09 lua1 = -6.118794686e-16
+ ub1 = -2.337858579e-18 lub1 = 8.983557464e-25 wub1 = -3.081487911e-39
+ uc1 = -8.386929930e-11 luc1 = 6.941675076e-17 wuc1 = 5.169878828e-32 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.42 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.215768093e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.945977550e-8
+ k1 = 3.667703539e-01 lk1 = 1.074781426e-7
+ k2 = 1.756159980e-02 lk2 = -3.063052309e-08 pk2 = -2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 7.575464332e-02 ldsub = 1.297992051e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.335627272e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.995746010e-9
+ nfactor = 2.533949421e+00 lnfactor = 1.593465777e-7
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 3.104053217e-02 lu0 = -4.183302695e-9
+ ua = -1.085244136e-09 lua = -2.610652142e-16
+ ub = 1.941064728e-18 lub = 8.127793964e-26
+ uc = 7.725809959e-11 luc = -7.422229282e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.854301274e+04 lvsat = 2.656444100e-2
+ a0 = 1.5
+ ags = 2.399526108e+00 lags = -6.206694043e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.102885254e-02 lketa = -2.318523268e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.820641385e-01 lpclm = -4.191721304e-8
+ pdiblc1 = 8.594644286e-01 lpdiblc1 = -1.836093976e-7
+ pdiblc2 = -4.584242403e-04 lpdiblc2 = 7.927530709e-10
+ pdiblcb = 1.836288000e-01 lpdiblcb = -1.065646702e-07 wpdiblcb = 1.110223025e-22 ppdiblcb = -5.551115123e-29
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.177411360e-06 lalpha0 = 3.196940107e-14
+ alpha1 = 0.85
+ beta0 = 1.686115330e+01 lbeta0 = 5.909010965e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.134635824e-01 lkt1 = 1.750969425e-8
+ kt2 = -5.758888667e-02 lkt2 = 1.055600904e-8
+ at = 7.152581445e+04 lat = -1.273506899e-2
+ ute = -2.267519941e+00 lute = 5.181754085e-7
+ ua1 = -3.630814747e-10 lua1 = 7.175291234e-16
+ ub1 = 3.233485706e-19 lub1 = -4.609516086e-25 pub1 = -3.851859889e-46
+ uc1 = 5.335421127e-11 luc1 = -6.750973096e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.43 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {7.248237971e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.638514448e-08 wvth0 = -2.394712385e-07 pvth0 = 6.245074640e-14
+ k1 = 4.295684749e-01 lk1 = 9.110127180e-8
+ k2 = 1.435086712e-01 lk2 = -6.347575604e-08 wk2 = -1.533740585e-07 pk2 = 3.999780722e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.865102111e-01 ldsub = -8.163449643e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 1.452502183e-02 lcdscd = -2.379677943e-9
+ cit = 0.0
+ voff = {2.523976002e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.440921144e-8
+ nfactor = -1.535733464e+00 lnfactor = 1.220662899e-06 wnfactor = 1.453221104e-05 pnfactor = -3.789797188e-12
+ eta0 = 1.823610115e+00 leta0 = -3.477868474e-7
+ etab = 1.175887311e-01 letab = -3.082848608e-08 petab = -4.336808690e-30
+ u0 = -5.000498844e-02 lu0 = 1.695223444e-08 wu0 = 4.063791962e-08 pu0 = -1.059780050e-14
+ ua = -4.324870790e-09 lua = 5.837840623e-16 wua = -6.692985545e-16 pua = 1.745436928e-22
+ ub = 1.603646406e-18 lub = 1.692719142e-25 wub = 3.889697840e-24 pub = -1.014378741e-30
+ uc = -1.902958301e-10 luc = 6.903209619e-17 wuc = 4.594129313e-16 puc = -1.198084607e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.974749511e+05 lvsat = -1.843483487e-03 wvsat = -9.136585120e-02 pvsat = 2.382693487e-8
+ a0 = 1.5
+ ags = -3.334129838e+00 lags = 8.745877952e-07 wags = 1.554312234e-21 pags = -8.326672685e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.455082892e-01 lketa = 1.057719111e-07 wketa = 4.665307035e-07 pketa = -1.216646760e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.154275872e-01 lpclm = -7.669653339e-08 wpclm = 3.105476395e-07 ppclm = -8.098647672e-14
+ pdiblc1 = -3.939770822e-01 lpdiblc1 = 1.432706002e-7
+ pdiblc2 = -1.329380080e-02 lpdiblc2 = 4.140039583e-09 ppdiblc2 = 3.469446952e-30
+ pdiblcb = -5.567066175e-01 lpdiblcb = 8.650444195e-8
+ drout = 2.353690284e+00 ldrout = -3.530234743e-7
+ pscbe1 = 8.233852396e+08 lpscbe1 = -6.098543103e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.221243171e-05 lalpha0 = -2.324237417e-12
+ alpha1 = 0.85
+ beta0 = 3.294674335e+01 lbeta0 = -3.603995590e-06 wbeta0 = 1.013206002e-06 pbeta0 = -2.642299403e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 6.837569132e-03 lkt1 = -6.602036187e-08 wkt1 = -5.066030008e-07 pkt1 = 1.321149702e-13
+ kt2 = 1.496186997e-02 lkt2 = -8.364212580e-9
+ at = -8.095366830e+04 lat = 2.702944539e-2
+ ute = 2.549898990e+00 lute = -7.381400046e-7
+ ua1 = 8.962747083e-09 lua1 = -1.714516403e-15
+ ub1 = -7.309374636e-18 lub1 = 1.529555746e-24
+ uc1 = -2.120305980e-10 luc1 = 6.853354557e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.44 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.816972340e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 8.786277135e-8
+ k1 = 0.90707349
+ k2 = -1.891979008e-01 wk2 = 5.627343775e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 4.862340286e+00 wnfactor = -5.331915197e-6
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 3.884972020e-02 wu0 = -1.491018404e-8
+ ua = -1.264981373e-09 wua = 2.455678028e-16
+ ub = 2.490880869e-18 wub = -1.427142709e-24
+ uc = 1.715341584e-10 wuc = -1.685600893e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.878123790e+05 wvsat = 3.352242609e-2
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.088925112e-01 wketa = -1.711716229e-7
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.134246447e-01 wpclm = -1.139409326e-7
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.405649150e+01 wbeta0 = -3.717485566e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.392064900e-01 wkt1 = 1.858742783e-7
+ kt2 = -0.028878939
+ at = 60720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.45 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.171504489e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.631718124e-07 wvth0 = 4.720315981e-09 pvth0 = 3.296096131e-13
+ k1 = 4.555796457e-01 lk1 = 6.197035863e-06 wk1 = 1.329169773e-07 pk1 = -9.384885502e-12
+ k2 = 6.474164105e-03 lk2 = -2.592850776e-06 wk2 = -5.341824451e-08 pk2 = 3.948676993e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.018345153e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.328226721e-07 wvoff = -2.874894333e-09 pvoff = -4.315619939e-13
+ nfactor = 3.068193461e+00 lnfactor = -5.376638958e-05 wnfactor = -9.389192773e-07 pnfactor = 8.357530486e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.091953141e-02 lu0 = 1.864391935e-07 wu0 = 1.118635428e-09 pu0 = -3.112530291e-13
+ ua = -7.558861509e-10 lua = -1.482132562e-15 wua = 4.467832666e-17 pua = 3.012020984e-21
+ ub = 1.549535476e-18 lub = 1.380658775e-23 wub = -2.760243305e-26 pub = -2.415799785e-29
+ uc = -7.319592212e-11 luc = 5.364165217e-15 wuc = 1.790877147e-16 puc = -7.480901143e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.090524119e+00 la0 = 1.129571087e-05 wa0 = 4.310059281e-07 pa0 = -1.521223700e-11
+ ags = 3.090914179e-01 lags = 4.137844151e-06 wags = 1.099036507e-07 pags = -6.054113547e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.198190121e-24 lb0 = 3.418877166e-28 wb0 = 1.363034970e-29 pb0 = -4.545573362e-34
+ b1 = 0.0
+ keta = -5.303646030e-03 lketa = -2.334581660e-07 wketa = -1.596515128e-09 pketa = 3.877846151e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.242116906e-02 lpclm = 6.225321695e-07 wpclm = 3.583640978e-08 ppclm = -7.171147271e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 6.355388330e-03 lpdiblc2 = -1.156498144e-07 wpdiblc2 = -4.682491401e-09 ppdiblc2 = 1.530420327e-13
+ pdiblcb = 9.324003944e+00 lpdiblcb = -2.529245211e-04 wpdiblcb = -1.371827341e-05 ppdiblcb = 2.997970971e-10
+ drout = 0.56
+ pscbe1 = 3.084204719e+08 lpscbe1 = 1.146351867e+04 wpscbe1 = 5.680178049e+02 ppscbe1 = -1.412739309e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.376827215e-01 lkt1 = -8.824353779e-07 wkt1 = 1.771038384e-08 pkt1 = 1.704077709e-12
+ kt2 = -4.786010220e-02 lkt2 = -9.849535387e-07 wkt2 = 1.946113545e-09 pkt2 = 1.723185705e-12
+ at = 140000.0
+ ute = -1.882501289e+00 lute = -2.573942053e-05 wute = -3.860869844e-08 pute = 4.413345560e-11
+ ua1 = 6.966609528e-10 lua1 = -6.345000468e-14 wua1 = -7.160395961e-16 pua1 = 1.025617504e-19
+ ub1 = -1.119883260e-18 lub1 = 4.227123315e-23 wub1 = 9.492126458e-25 pub1 = -6.358906180e-29
+ uc1 = -3.282482510e-12 luc1 = 2.541245255e-15 wuc1 = 3.265619405e-17 puc1 = -4.067790957e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.46 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.089962558e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.119191350e-8
+ k1 = 7.652644259e-01 wk1 = -3.360743707e-7
+ k2 = -1.230984961e-01 wk2 = 1.439091864e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.019965643e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -2.444136323e-8
+ nfactor = 3.813230110e-01 wnfactor = 3.237593572e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 4.023646647e-02 wu0 = -1.443562762e-8
+ ua = -8.299528348e-10 wua = 1.951982005e-16
+ ub = 2.239492770e-18 wub = -1.234851256e-24
+ uc = 1.948677720e-10 wuc = -1.947557287e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.655005238e+00 wa0 = -3.291959449e-7
+ ags = 5.158721086e-01 wags = -1.926388654e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.886981675e-24 wb0 = -9.085266575e-30
+ b1 = 0.0
+ keta = -1.697026253e-02 wketa = 1.778226465e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 5.760144238e-04 wpdiblc2 = 2.965485678e-9
+ pdiblcb = -3.315405677e+00 wpdiblcb = 1.263501771e-6
+ drout = 0.56
+ pscbe1 = 8.812874582e+08 wpscbe1 = -1.379711096e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.817807084e-01 wkt1 = 1.028683436e-7
+ kt2 = -9.708123418e-02 wkt2 = 8.805895814e-8
+ at = 140000.0
+ ute = -3.168778627e+00 wute = 2.166874665e-6
+ ua1 = -2.474129274e-09 wua1 = 4.409283838e-15
+ ub1 = 9.925391686e-19 wub1 = -2.228526689e-24
+ uc1 = 1.237112925e-10 wuc1 = -1.706237249e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.47 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.910522174e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.437458519e-07 wvth0 = 2.997572762e-08 pvth0 = -7.036525518e-14
+ k1 = 7.994523375e-01 lk1 = -2.738720441e-07 wk1 = -3.947886715e-07 pk1 = 4.703476985e-13
+ k2 = -1.351107206e-01 lk2 = 9.622735951e-08 wk2 = 1.684724982e-07 pk2 = -1.967714338e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.299661719e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.770200590e-08 wvoff = -3.898426245e-08 pvoff = 1.165000535e-13
+ nfactor = 1.858059204e-01 lnfactor = 1.566245571e-06 wnfactor = 3.782761542e-06 pnfactor = -4.367223944e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.891653727e-02 lu0 = 1.057367036e-08 wu0 = -1.244101576e-08 pu0 = -1.597840875e-14
+ ua = -9.813544586e-10 lua = 1.212846008e-15 wua = 4.137751516e-16 pua = -1.750973179e-21
+ ub = 2.304602062e-18 lub = -5.215766049e-25 wub = -1.321137456e-24 pub = 6.912202832e-31
+ uc = 2.324585165e-10 luc = -3.011314097e-16 wuc = -2.375702840e-16 puc = 3.429782407e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.513699368e+00 la0 = 1.131971079e-06 wa0 = -1.427725248e-08 pa0 = -2.522746252e-12
+ ags = 3.813023510e-01 lags = 1.078009531e-06 wags = -2.665599029e-08 pags = -1.329653292e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.579523060e-23 lb0 = -6.335128974e-29 wb0 = -1.819503157e-29 pb0 = 7.297637790e-35
+ b1 = 0.0
+ keta = -4.569511354e-03 lketa = -9.933976387e-08 wketa = -9.546900219e-09 pketa = 2.189280913e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.010244142e-01 lpclm = 2.279512528e-06 wpclm = -1.915501765e-07 ppclm = 1.534467472e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.750100865e-03 lpdiblc2 = 2.664479779e-08 wpdiblc2 = 6.572556201e-09 ppdiblc2 = -2.889547005e-14
+ pdiblcb = -6.614683933e+00 lpdiblcb = 2.642981206e-05 wpdiblcb = 2.530410575e-06 ppdiblcb = -1.014893531e-11
+ drout = 0.56
+ pscbe1 = 8.121675033e+08 lpscbe1 = 5.537051663e+02 wpscbe1 = -3.953947846e+01 ppscbe1 = -7.885147326e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.768321321e-01 lkt1 = -3.964198524e-08 wkt1 = 9.858861725e-08 pkt1 = 3.428397196e-14
+ kt2 = -9.312253560e-02 lkt2 = -3.171228714e-08 wkt2 = 8.357010014e-08 pkt2 = 3.595928076e-14
+ at = 140000.0
+ ute = -2.715161340e+00 lute = -3.633831010e-06 wute = 1.410789675e-06 pute = 6.056835047e-12
+ ua1 = -2.027849365e-09 lua1 = -3.575052845e-15 wua1 = 3.777501339e-15 pua1 = 5.061074396e-21
+ ub1 = 6.961711965e-19 lub1 = 2.374140402e-24 wub1 = -1.879958151e-24 pub1 = -2.792307964e-30
+ uc1 = 9.557869579e-11 luc1 = 2.253642120e-16 wuc1 = -1.452897767e-16 puc1 = -2.029448378e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.48 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.078368527e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.246523284e-07 wvth0 = -1.120050086e-07 pvth0 = 4.990890939e-13
+ k1 = 8.120910460e-01 lk1 = -3.245631992e-07 wk1 = -4.276800911e-07 pk1 = 6.022681437e-13
+ k2 = -1.644818103e-01 lk2 = 2.140285150e-07 wk2 = 2.109338787e-07 pk2 = -3.670749443e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.625454835e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.613514734e-07 wvoff = 8.810008177e-08 pvoff = -3.932080551e-13
+ nfactor = -2.962307874e+00 lnfactor = 1.419265630e-05 wnfactor = 7.501482573e-06 pnfactor = -1.928221819e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 4.471392842e-02 lu0 = -1.267842493e-08 wu0 = -1.771484690e-08 pu0 = 5.173799349e-15
+ ua = -1.553357880e-09 lua = 3.507029322e-15 wua = 1.511181270e-15 pua = -6.152434275e-21
+ ub = 3.913268596e-18 lub = -6.973593817e-24 wub = -3.748765726e-24 pub = 1.042791776e-29
+ uc = 2.235302459e-10 luc = -2.653220272e-16 wuc = -2.615174968e-16 puc = 4.390253863e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 3.535560920e-01 la0 = 5.785057490e-06 wa0 = 1.338507215e-06 pa0 = -7.948475256e-12
+ ags = 4.463057386e-01 lags = 8.172948537e-07 wags = -3.567002700e-07 pags = -5.916316050e-15
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.929516167e-24 lb0 = 3.180359243e-29 wb0 = 9.134263418e-30 pb0 = -3.663557584e-35
+ b1 = 0.0
+ keta = -8.468260840e-02 lketa = 2.219767242e-07 wketa = 1.303367018e-07 pketa = -3.421151014e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.760744296e-01 lpclm = -3.510743488e-08 wpclm = 1.532375006e-07 ppclm = 1.515978842e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 4.167704910e-03 lpdiblc2 = -1.101040765e-09 wpdiblc2 = -3.209128685e-09 ppdiblc2 = 1.033677475e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.132630470e+09 lpscbe1 = -7.316032133e+02 wpscbe1 = -5.096940303e+02 ppscbe1 = 1.097174562e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.677224275e-01 lkt1 = -7.617906097e-08 wkt1 = 8.290625060e-08 pkt1 = 9.718258858e-14
+ kt2 = -9.481774513e-02 lkt2 = -2.491316450e-08 wkt2 = 8.190650560e-08 pkt2 = 4.263160247e-14
+ at = 1.542800880e+05 lat = -5.727437697e-02 wat = 1.690486752e-02 pat = -6.780180599e-8
+ ute = -2.460414528e+00 lute = -4.655565958e-06 wute = 8.159235804e-07 pute = 8.442715652e-12
+ ua1 = 2.043774588e-09 lua1 = -1.990546520e-14 wua1 = -3.173685068e-15 pua1 = 3.294079552e-20
+ ub1 = -3.427478360e-18 lub1 = 1.891321631e-23 wub1 = 4.926560507e-24 pub1 = -3.009179771e-29
+ uc1 = 5.219392052e-11 luc1 = 3.993712613e-16 wuc1 = -6.736468393e-17 puc1 = -5.154857089e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.49 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {3.607891851e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.721076630e-07 wvth0 = 1.997891469e-07 pvth0 = -1.278622288e-13
+ k1 = 7.207257604e-01 lk1 = -1.408471619e-07 wk1 = -1.388077264e-07 pk1 = 2.140763709e-14
+ k2 = -7.661043593e-02 lk2 = 3.733798554e-08 wk2 = 2.904935389e-08 pk2 = -1.344088184e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {2.102585095e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.077711959e-07 wvoff = -1.395073933e-07 pvoff = 6.446186923e-14
+ nfactor = 4.244063249e+00 lnfactor = -2.978138602e-07 wnfactor = -1.710079880e-06 pnfactor = -7.597373725e-13
+ eta0 = 1.583044666e-01 leta0 = -1.574535251e-07 weta0 = -2.178916211e-13 peta0 = 4.381334211e-19
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 4.680736892e-02 lu0 = -1.688788579e-08 wu0 = -2.180686675e-08 pu0 = 1.340197559e-14
+ ua = 2.141002321e-09 lua = -3.921538449e-15 wua = -3.523531124e-15 pua = 3.971294921e-21
+ ub = -1.868587428e-18 lub = 4.652481330e-24 wub = 3.881027802e-24 pub = -4.913964248e-30
+ uc = 9.535499624e-11 luc = -7.589029566e-18 wuc = -6.621778757e-17 puc = 4.631946528e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.244250068e+05 lvsat = -8.932918177e-02 wvsat = -6.281815435e-02 pvsat = 1.263138653e-7
+ a0 = 4.283641088e+00 la0 = -2.117502399e-06 wa0 = -3.287048110e-06 pa0 = 1.352526634e-12
+ ags = -1.023502674e+00 lags = 3.772765031e-06 wags = 1.600763217e-06 pags = -3.941956491e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.585903233e-23 lb0 = -1.603008786e-29 wb0 = -1.826852684e-29 pb0 = 1.846557117e-35
+ b1 = 0.0
+ keta = 2.722724700e-01 lketa = -4.957835501e-07 wketa = -3.452300349e-07 pketa = 6.141478349e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.346917266e-01 lpclm = 2.198405601e-06 wpclm = 1.335257817e-06 ppclm = -2.225192019e-12
+ pdiblc1 = -6.244660677e-01 lpdiblc1 = 2.039874166e-06 wpdiblc1 = 1.228322048e-06 ppdiblc1 = -2.469892777e-12
+ pdiblc2 = 1.096863474e-02 lpdiblc2 = -1.477625526e-08 wpdiblc2 = -7.126979603e-09 ppdiblc2 = 1.821473452e-14
+ pdiblcb = -1.864189408e-01 lpdiblcb = 3.245789463e-07 wpdiblcb = 2.143219745e-07 ppdiblcb = -4.309556259e-13
+ drout = 1.243869036e+00 ldrout = -1.375114283e-06 wdrout = -5.983295634e-07 pdrout = 1.203112709e-12
+ pscbe1 = 2.175922303e+09 lpscbe1 = -2.829439825e+03 wpscbe1 = -1.584968930e+03 ppscbe1 = 3.259322276e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.227897527e-08 lalpha0 = 2.257689916e-13 walpha0 = 1.307349726e-13 palpha0 = -2.628800527e-19
+ alpha1 = -4.102156589e-01 lalpha1 = 2.534024004e-06 walpha1 = 1.629829325e-06 palpha1 = -3.277237990e-12
+ beta0 = 1.132913022e+01 lbeta0 = 5.089037525e-06 wbeta0 = 2.915389890e-06 pbeta0 = -5.862225174e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.625754292e-01 lkt1 = 3.156286268e-07 wkt1 = 2.712540534e-07 pkt1 = -2.815445364e-13
+ kt2 = -1.804497844e-01 lkt2 = 1.472745412e-07 wkt2 = 2.090513359e-07 pkt2 = -2.130294423e-13
+ at = 2.422931815e+05 lat = -2.342498731e-01 wat = -1.213367992e-01 pat = 2.101726021e-7
+ ute = -8.065528057e+00 lute = 6.615117856e-06 wute = 9.531225997e-06 pute = -9.081892433e-12
+ ua1 = -1.852321893e-08 lua1 = 2.145035744e-14 wua1 = 2.824977458e-14 pua1 = -3.024505721e-20
+ ub1 = 1.537495432e-17 lub1 = -1.889445208e-23 wub1 = -2.315483117e-23 pub1 = 2.637387153e-29
+ uc1 = 6.118300250e-10 luc1 = -7.259371827e-16 wuc1 = -7.957964577e-16 puc1 = 9.492347038e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.50 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.006127632e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.077594773e-08 wvth0 = 1.118488580e-07 pvth0 = -3.897341593e-14
+ k1 = 5.472829464e-01 lk1 = 3.446640629e-08 wk1 = -1.774588569e-07 pk1 = 6.047565865e-14
+ k2 = -2.083649143e-02 lk2 = -1.903753673e-08 wk2 = 3.082269978e-08 pk2 = -3.136561385e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.423481142e-01 ldsub = 1.189208791e-07 wdsub = 7.273859612e-08 pdsub = -7.352315462e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-4.744689245e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.855990548e-08 wvoff = -1.266209824e-07 pvoff = 5.143646549e-14
+ nfactor = 5.440351800e+00 lnfactor = -1.507005579e-06 wnfactor = -5.548086719e-06 pnfactor = 3.119666208e-12
+ eta0 = -4.954534531e-01 leta0 = 5.033558275e-07 weta0 = 4.357832419e-13 peta0 = -2.225919791e-19
+ etab = -1.690560735e-01 letab = 8.559444360e-08 wetab = -1.376354510e-09 petab = 1.391199869e-15
+ u0 = 3.385321651e-02 lu0 = -3.794009886e-09 wu0 = -1.153959056e-08 pu0 = 3.023956554e-15
+ ua = -1.573012728e-09 lua = -1.674640342e-16 wua = 3.305082081e-16 pua = 7.568592061e-23
+ ub = 2.487104708e-18 lub = 2.498086988e-25 wub = -5.754597958e-25 pub = -4.094089753e-31
+ uc = 1.050098941e-10 luc = -1.734806517e-17 wuc = -4.886661494e-17 puc = 2.878114290e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.943727398e+04 lvsat = 8.640837759e-02 wvsat = 9.220300603e-02 pvsat = -3.037935331e-8
+ a0 = 2.892326084e+00 la0 = -7.111806710e-07 wa0 = -3.939951154e-06 pa0 = 2.012471890e-12
+ ags = 4.016569868e+00 lags = -1.321669733e-06 wags = -4.254988253e-06 pags = 1.976955114e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.938196835e-01 lketa = 1.774930733e-07 wketa = 5.131068521e-07 pketa = -2.534470738e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.783136245e+00 lpclm = -1.357365663e-06 wpclm = -2.191497666e-06 ppclm = 1.339603049e-12
+ pdiblc1 = 1.303826661e+00 lpdiblc1 = 9.078287259e-08 wpdiblc1 = -8.804167052e-07 ppdiblc1 = -3.384091679e-13
+ pdiblc2 = -7.060664760e-03 lpdiblc2 = 3.447508269e-09 wpdiblc2 = 1.976580268e-08 ppdiblc2 = -8.968113309e-15
+ pdiblcb = 2.978378816e-01 lpdiblcb = -1.649010702e-07 wpdiblcb = -4.286439490e-07 ppdiblcb = 2.189453282e-13
+ drout = -1.257229751e+00 ldrout = 1.152961356e-06 wdrout = 1.196659127e-06 pdrout = -6.112367287e-13
+ pscbe1 = -2.077353648e+09 lpscbe1 = 1.469711960e+03 wpscbe1 = 3.314515743e+03 ppscbe1 = -1.693008238e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.201866089e-05 lalpha0 = 1.229089672e-11 walpha0 = 1.387644358e-11 palpha0 = -1.415684987e-17
+ alpha1 = 3.370431318e+00 lalpha1 = -1.287401031e-06 walpha1 = -3.259658651e-06 palpha1 = 1.664988004e-12
+ beta0 = 3.023906564e+00 lbeta0 = 1.348384132e-05 wbeta0 = 1.248244278e-05 pbeta0 = -1.553246830e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.972282506e-01 lkt1 = -5.365918644e-08 wkt1 = -5.181921065e-08 pkt1 = 4.501339586e-14
+ kt2 = -3.092003953e-02 lkt2 = -3.868031485e-09 wkt2 = -5.967831825e-09 pkt2 = 4.308922176e-15
+ at = -1.637544366e+04 lat = 2.720875177e-02 wat = 1.594765612e-01 pat = -7.366961124e-8
+ ute = -1.718773352e+00 lute = 1.999070543e-07 wute = 9.848824781e-07 pute = -4.433680528e-13
+ ua1 = 4.536080362e-09 lua1 = -1.857659456e-15 wua1 = -3.609925333e-15 pua1 = 1.958281428e-21
+ ub1 = -6.397761641e-18 lub1 = 3.113104392e-24 wub1 = 6.381891540e-24 pub1 = -3.481434268e-30
+ uc1 = -3.041207366e-10 luc1 = 1.998930238e-16 wuc1 = 3.462202823e-16 puc1 = -2.050998288e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.51 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.086461845e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.440601139e-08 wvth0 = 2.032606287e-08 pvth0 = 7.775146479e-15
+ k1 = 8.102388335e-01 lk1 = -9.984777950e-08 wk1 = -6.971022941e-07 pk1 = 3.259022514e-13
+ k2 = -1.499352824e-01 lk2 = 4.690431832e-08 wk2 = 2.632937091e-07 pk2 = -1.218794983e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.602808753e-01 ldsub = 2.734995301e-07 wdsub = 3.710317849e-07 pdsub = -2.258871393e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = -4.178715321e-03 lcdscd = 4.892673684e-09 wcdscd = 1.505708913e-08 pcdscd = -7.690950329e-15
+ cit = 0.0
+ voff = {-1.955161298e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.707178801e-08 wvoff = 9.738653616e-08 pvoff = -6.298343888e-14
+ nfactor = -2.910502403e+00 lnfactor = 2.758493836e-06 wnfactor = 8.558308045e-06 pnfactor = -4.085682748e-12
+ eta0 = -9.099168273e-01 leta0 = 7.150579165e-07 weta0 = 2.200574058e-06 peta0 = -1.124022421e-12
+ etab = -1.264674471e-01 letab = 6.384076948e-08 wetab = 1.978157696e-07 petab = -1.003533484e-13
+ u0 = 4.874596896e-02 lu0 = -1.140101934e-08 wu0 = -2.783174266e-08 pu0 = 1.134575976e-14
+ ua = 1.098853166e-09 lua = -1.532215726e-15 wua = -3.433252440e-15 pua = 1.998162167e-21
+ ub = 1.624399029e-19 lub = 1.437214936e-24 wub = 2.795877278e-24 pub = -2.131440754e-30
+ uc = 1.194575444e-10 luc = -2.472772268e-17 wuc = -6.633465772e-17 puc = 3.770357460e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.239741596e+04 lvsat = 1.906906366e-02 wvsat = 9.660460239e-03 pvsat = 1.178222349e-8
+ a0 = 1.5
+ ags = 6.419781951e+00 lags = -2.549196820e-06 wags = -6.319568808e-06 pags = 3.031513958e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.766946049e-01 lketa = 6.658862296e-08 wketa = 2.289766575e-07 pketa = -1.083173482e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.150865120e-01 lpclm = 2.251631461e-07 wpclm = 1.253066616e-06 ppclm = -4.198321631e-13
+ pdiblc1 = 3.441624505e+00 lpdiblc1 = -1.001174337e-06 wpdiblc1 = -4.058980054e-06 ppdiblc1 = 1.285156491e-12
+ pdiblc2 = 1.333581783e-02 lpdiblc2 = -6.970729485e-09 wpdiblc2 = -2.168361052e-08 ppdiblc2 = 1.220366666e-14
+ pdiblcb = 5.318277763e-01 lpdiblcb = -2.844198325e-07 wpdiblcb = -5.473451131e-07 ppdiblcb = 2.795762210e-13
+ drout = -4.209953797e-01 ldrout = 7.258245460e-07 wdrout = 2.233708109e-06 pdrout = -1.140946830e-12
+ pscbe1 = 7.754520529e+08 lpscbe1 = 1.253874771e+01 wpscbe1 = 3.858770358e+01 ppscbe1 = -1.971005876e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.178576889e-05 lalpha0 = 1.319272505e-13 walpha0 = -1.353175267e-11 palpha0 = -1.571269422e-19
+ alpha1 = 0.85
+ beta0 = 2.640847418e+01 lbeta0 = 1.539331569e-06 wbeta0 = -1.500773919e-05 pbeta0 = -1.490868209e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.453160813e-01 lkt1 = 2.198200426e-08 wkt1 = 5.006996227e-08 pkt1 = -7.030167216e-15
+ kt2 = -9.446450759e-02 lkt2 = 2.858959318e-08 wkt2 = 5.796596854e-08 pkt2 = -2.834756798e-14
+ at = 6.895266352e+04 lat = -1.637565078e-02 wat = 4.044818287e-03 pat = 5.722747009e-9
+ ute = -5.390597267e+00 lute = 2.075423305e-06 wute = 4.909265188e-06 pute = -2.447887800e-12
+ ua1 = -7.555439804e-09 lua1 = 4.318519763e-15 wua1 = 1.130589821e-14 pua1 = -5.660512418e-21
+ ub1 = 7.044167282e-18 lub1 = -3.752844715e-24 wub1 = -1.056467000e-23 pub1 = 5.174632115e-30
+ uc1 = 4.011161556e-10 luc1 = -1.603321074e-16 wuc1 = -5.466581287e-16 puc1 = 2.509699632e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.52 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.009440125e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.681207239e-09 wvth0 = 1.124525592e-07 pvth0 = -1.625015399e-14
+ k1 = -8.800822560e-01 lk1 = 3.409642962e-07 wk1 = 2.058681893e-06 pk1 = -3.927676836e-13
+ k2 = 5.270626092e-01 lk2 = -1.296472538e-07 wk2 = -7.562947674e-07 pk2 = 1.440149021e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.060018301e+00 ldsub = -3.055234108e-07 wdsub = -1.844674918e-06 pdsub = 3.519381490e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.873471940e-02 lcdscd = -8.906409304e-09 wcdscd = -5.377531833e-08 pcdscd = 1.025957788e-14
+ cit = 0.0
+ voff = {3.668248164e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.095788580e-07 wvoff = -5.369484809e-07 pvoff = 1.024422529e-13
+ nfactor = 2.625586680e+01 lnfactor = -4.847686923e-06 wnfactor = -2.915429475e-05 pnfactor = 5.749236084e-12
+ eta0 = 6.823313069e+00 leta0 = -1.301660175e-06 weta0 = -7.859193065e-06 peta0 = 1.499424008e-12
+ etab = 5.607718891e-01 letab = -1.153816281e-07 wetab = -6.966537879e-07 petab = 1.329117896e-13
+ u0 = -6.200883872e-02 lu0 = 1.748228394e-08 wu0 = 5.950715600e-08 pu0 = -1.143100227e-14
+ ua = -1.466912303e-08 lua = 2.579851715e-15 wua = 1.559116256e-14 pua = -2.963138924e-21
+ ub = 1.883521419e-17 lub = -3.432383179e-24 wub = -2.319715496e-23 pub = 4.647178152e-30
+ uc = 4.150765126e-11 luc = -4.399481842e-18 wuc = 9.503362116e-17 puc = -4.379013379e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.049693872e+05 lvsat = -1.289599042e-02 wvsat = -1.031465950e-01 pvsat = 4.120072420e-8
+ a0 = 1.5
+ ags = -1.590700091e+01 lags = 3.273315576e-06 wags = 1.976369838e-05 pags = -3.770636959e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.929877674e-01 lketa = -5.589796420e-08 wketa = -6.943348799e-07 pketa = 1.324693744e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.658623088e+00 lpclm = -2.895526856e-07 wpclm = -1.329284751e-06 ppclm = 2.536089204e-13
+ pdiblc1 = -2.453601965e+00 lpdiblc1 = 5.362181932e-07 wpdiblc1 = 3.237590262e-06 ppdiblc1 = -6.176868957e-13
+ pdiblc2 = -7.281004859e-02 lpdiblc2 = 1.549490643e-08 wpdiblc2 = 9.355549441e-08 ppdiblc2 = -1.784907856e-14
+ pdiblcb = -1.800274390e+00 lpdiblcb = 3.237597630e-07 wpdiblcb = 1.954803975e-06 ppdiblcb = -3.729492313e-13
+ drout = 7.428673782e+00 ldrout = -1.321259276e-06 wdrout = -7.977528961e-06 pdrout = 1.522000840e-12
+ pscbe1 = 9.110564793e+08 lpscbe1 = -2.282498823e+01 wpscbe1 = -1.378132271e+02 ppscbe1 = 2.629283434e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 4.571095995e-05 lalpha0 = -8.715287625e-12 walpha0 = -5.265740848e-11 palpha0 = 1.004629633e-17
+ alpha1 = 0.85
+ beta0 = 8.293324901e+01 lbeta0 = -1.320153836e-05 wbeta0 = -7.756218182e-05 pbeta0 = 1.482245466e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.702197084e-01 lkt1 = 2.847652154e-08 wkt1 = 8.610539949e-08 pkt1 = -1.642770475e-14
+ kt2 = 1.352038480e-01 lkt2 = -3.130469859e-08 wkt2 = -1.890122130e-07 pkt2 = 3.606088406e-14
+ at = -2.920533911e+05 lat = 7.776967419e-02 wat = 3.318344095e-01 pat = -7.976018933e-8
+ ute = 1.316122831e+01 lute = -2.762633080e-06 wute = -1.668028812e-05 pute = 3.182365449e-12
+ ua1 = 3.361023680e-08 lua1 = -6.416912376e-15 wua1 = -3.874417781e-14 pua1 = 7.391846708e-21
+ ub1 = -2.929791289e-17 lub1 = 5.724661006e-24 wub1 = 3.456448692e-23 pub1 = -6.594420202e-30
+ uc1 = -1.197252937e-09 luc1 = 2.565001747e-16 wuc1 = 1.548702521e-15 puc1 = -2.954707592e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.53 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.202389672e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.727778751e-8
+ k1 = 0.90707349
+ k2 = -1.524801971e-01 wk2 = -1.444295688e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 8.468382376e-01 wnfactor = 9.801809689e-7
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 2.962411096e-02 wu0 = -4.081536500e-10
+ ua = -1.146895435e-09 wua = 5.994473803e-17
+ ub = 8.444644532e-19 wub = 1.160911940e-24
+ uc = 1.844787831e-11 wuc = 7.208113314e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.373753791e+05 wvsat = 1.128059602e-1
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 0.0
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.14094
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.373771914e+01 wbeta0 = 1.293399123e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.22096074
+ kt2 = -0.028878939
+ at = 1.155743918e+05 wat = -8.622660822e-2
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.54 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.984260027e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.422502814e-06 wvth0 = -2.040967952e-07 pvth0 = 4.084137293e-12
+ k1 = 5.000310512e-01 lk1 = -5.305874165e-07 wk1 = 8.171198085e-08 pk1 = -1.635120962e-12
+ k2 = -3.823891573e-02 lk2 = 8.018114364e-07 wk2 = -1.911817029e-09 pk2 = 3.825696143e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.348192401e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.589023715e-07 wvoff = -1.249651158e-08 pvoff = 2.500650189e-13
+ nfactor = -4.099373251e+00 lnfactor = 1.459041087e-04 wnfactor = 7.317630180e-06 pnfactor = -1.464315316e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 7.069728418e-02 lu0 = -8.603134005e-07 wu0 = -4.470263087e-08 pu0 = 8.945347799e-13
+ ua = 7.554738052e-10 lua = -2.833474780e-14 wua = -1.696305570e-15 pua = 3.394440776e-20
+ ub = 2.407223415e-18 lub = -2.480763985e-23 wub = -1.015600616e-24 pub = 2.032296659e-29
+ uc = 1.784860171e-10 luc = -3.055387225e-15 wuc = -1.108327650e-16 puc = 2.217850741e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.820568239e+00 la0 = -9.031672940e-06 wa0 = -4.099552559e-07 pa0 = 8.203526896e-12
+ ags = 6.122520352e-01 lags = -5.275064012e-06 wags = -2.393167654e-07 pags = 4.788916579e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.134409340e-08 lb0 = -1.227543525e-12 wb0 = -7.066422420e-14 pb0 = 1.414046668e-18
+ b1 = -5.307138953e-08 lb1 = 1.062000219e-12 wb1 = 6.113463188e-14 pb1 = -1.223352036e-18
+ keta = -1.145550966e-02 lketa = 1.985500596e-07 wketa = 5.490013447e-09 pketa = -1.098594842e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.693917305e-01 lpclm = -5.720297905e-06 wpclm = -3.292921230e-07 ppclm = 6.589394206e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 8.732858526e-03 lpdiblc2 = -1.117099292e-07 wpdiblc2 = -7.421175400e-09 ppdiblc2 = 1.485035528e-13
+ pdiblcb = -1.324901929e+01 lpdiblcb = 2.207283363e-04 wpdiblcb = 1.228431438e-05 ppdiblcb = -2.458187862e-10
+ drout = 0.56
+ pscbe1 = 3.239655734e+09 lpscbe1 = -4.958956792e+04 wpscbe1 = -2.808565893e+03 ppscbe1 = 5.620161106e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.507945870e-01 lkt1 = 3.167999322e-06 wkt1 = 1.480075613e-07 pkt1 = -2.961747636e-12
+ kt2 = -9.567707948e-02 lkt2 = 1.501617896e-06 wkt2 = 5.702801982e-08 pkt2 = -1.141175501e-12
+ at = -1.010089968e+04 lat = 3.003636982e+00 wat = 1.729060296e-01 pat = -3.459985556e-6
+ ute = -4.810391969e+00 lute = 7.049183513e-05 wute = 3.334122267e-06 pute = -6.671840719e-11
+ ua1 = -3.313444255e-09 lua1 = 9.339122385e-14 wua1 = 3.903328917e-15 pua1 = -7.810867964e-20
+ ub1 = 3.230221434e-19 lub1 = -2.531528804e-23 wub1 = -7.129162608e-25 pub1 = 1.426601473e-29
+ uc1 = -5.492017226e-11 luc1 = 6.105660860e-16 wuc1 = 9.213930127e-17 puc1 = -1.843779840e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.55 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.5273931+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47351598
+ k2 = 0.0018300469
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.11141737+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.1919
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0277048
+ ua = -6.6049995e-10
+ ub = 1.16751e-18
+ uc = 2.5799e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.369228
+ ags = 0.348641
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0015333577
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0031503727
+ pdiblcb = -2.2185512
+ drout = 0.56
+ pscbe1 = 761513800.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.29248
+ kt2 = -0.020636654
+ at = 140000.0
+ ute = -1.2877
+ ua1 = 1.3536e-9
+ ub1 = -9.4206e-19
+ uc1 = -2.4408323e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.56 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.170743503e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.266129549e-8
+ k1 = 4.567336080e-01 lk1 = 1.344399904e-7
+ k2 = 1.114140034e-02 lk2 = -7.459125980e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.168391204e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.343248247e-8
+ nfactor = 3.469646931e+00 lnfactor = -2.224971222e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.811640691e-02 lu0 = -3.297294898e-9
+ ua = -6.221534367e-10 lua = -3.071857119e-16
+ ub = 1.157713655e-18 lub = 7.847642182e-26
+ uc = 2.622213792e-11 luc = -3.389667350e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.501305188e+00 la0 = -1.058042092e-6
+ ags = 3.581621046e-01 lags = -7.627153156e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.285724033e-02 lketa = 9.071320047e-08 wketa = -1.734723476e-24 pketa = -2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.673104246e-01 lpclm = 3.611594172e-06 wpclm = 1.110223025e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 2.955579854e-03 lpdiblc2 = 1.560443807e-9
+ pdiblcb = -4.418017311e+00 lpdiblcb = 1.761945233e-5
+ drout = 0.56
+ pscbe1 = 7.778430133e+08 lpscbe1 = -1.308098334e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912466833e-01 lkt1 = -9.879836114e-9
+ kt2 = -2.057476356e-02 lkt2 = -4.957910604e-10
+ at = 140000.0
+ ute = -1.490445232e+00 lute = 1.624148668e-6
+ ua1 = 1.251425227e-09 lua1 = 8.185002439e-16
+ ub1 = -9.358332547e-19 lub1 = -4.988112379e-26
+ uc1 = -3.054834705e-11 luc1 = 4.918641870e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.57 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.106045433e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.086103068e-7
+ k1 = 4.408190516e-01 lk1 = 1.982698706e-7
+ k2 = 1.863132370e-02 lk2 = -1.046317395e-07 wk2 = 6.938893904e-24
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.606520361e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.999511228e-8
+ nfactor = 3.549780143e+00 lnfactor = -2.546368387e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.933554941e-02 lu0 = -8.187014548e-9
+ ua = -2.414911465e-10 lua = -1.833940696e-15
+ ub = 6.589395849e-19 lub = 2.078952480e-24
+ uc = -3.494870781e-12 luc = 1.157988951e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.515523305e+00 la0 = -1.115067914e-6
+ ags = 1.366518094e-01 lags = 8.121588595e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.846356849e-02 lketa = -7.501572108e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.091009455e-01 lpclm = 9.649571892e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.381838483e-03 lpdiblc2 = 7.872383663e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.901616173e+08 lpscbe1 = 2.208614822e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.957509478e-01 lkt1 = 8.185804823e-9
+ kt2 = -2.371415082e-02 lkt2 = 1.209561941e-8
+ at = 1.689553184e+05 lat = -1.161335857e-1
+ ute = -1.752105721e+00 lute = 2.673612892e-6
+ ua1 = -7.113229936e-10 lua1 = 8.690663327e-15 pua1 = 3.308722450e-36
+ ub1 = 8.493023065e-19 lub1 = -7.209677841e-24
+ uc1 = -6.285819551e-12 luc1 = -4.812538692e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.58 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.342275017e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.110959292e-8
+ k1 = 6.002258295e-01 lk1 = -1.222630466e-7
+ k2 = -5.139249434e-02 lk2 = 3.617117345e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.000814656e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.181140900e-8
+ nfactor = 2.759531280e+00 lnfactor = -9.573470380e-7
+ eta0 = 1.583042774e-01 leta0 = -1.574531447e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 2.787667965e-02 lu0 = -5.253539668e-9
+ ua = -9.177990006e-10 lua = -4.740303314e-16
+ ub = 1.500559190e-18 lub = 3.866355608e-25
+ uc = 3.787088470e-11 luc = 3.262121312e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.989214000e+04 lvsat = 2.032474338e-2
+ a0 = 1.430132279e+00 la0 = -9.433648340e-7
+ ags = 3.661307571e-01 lags = 3.507258042e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.742407017e-02 lketa = 3.736236032e-08 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.244546611e-01 lpclm = 2.667012826e-7
+ pdiblc1 = 4.418486520e-01 lpdiblc1 = -1.042565435e-7
+ pdiblc2 = 4.781655300e-03 lpdiblc2 = 1.036079606e-9
+ pdiblcb = -3.645777836e-04 lpdiblcb = -4.953656210e-8
+ drout = 7.244550742e-01 ldrout = -3.306839609e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.121294320e-08 lalpha0 = -2.438969205e-15 walpha0 = -2.646977960e-29
+ alpha1 = 1.004650258e+00 lalpha1 = -3.109685737e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.270979414e-01 lkt1 = 7.121790080e-8
+ kt2 = 1.029101439e-03 lkt2 = -3.765776583e-8
+ at = 1.369598812e+05 lat = -5.179760850e-2
+ ute = 2.085940234e-01 lute = -1.268934703e-6
+ ua1 = 6.000602418e-09 lua1 = -4.805582324e-15 wua1 = 3.308722450e-30
+ ub1 = -4.725912025e-18 lub1 = 4.000885084e-24
+ uc1 = -7.900628978e-11 luc1 = 9.809991654e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.59 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.977095171e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.057139584e-9
+ k1 = 3.932297063e-01 lk1 = 8.696573668e-8
+ k2 = 5.920903785e-03 lk2 = -2.176040699e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.054929839e-01 ldsub = 5.509492874e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.573674280e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.092439875e-9
+ nfactor = 6.240200030e-01 lnfactor = 1.201197864e-6
+ eta0 = -4.954530748e-01 leta0 = 5.033556343e-07 weta0 = -4.163336342e-23 peta0 = 1.058181320e-28
+ etab = -1.702508963e-01 letab = 8.680215367e-8
+ u0 = 2.383561950e-02 lu0 = -1.168892645e-9
+ ua = -1.286096305e-09 lua = -1.017605720e-16
+ ub = 1.987544147e-18 lub = -1.056020158e-25
+ uc = 6.258845349e-11 luc = 7.637040637e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.060478235e+04 lvsat = 6.003585447e-2
+ a0 = -5.279722970e-01 la0 = 1.035859858e-6
+ ags = 3.227856408e-01 lags = 3.945384409e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.161186290e-02 lketa = -4.252605433e-08 wketa = -1.387778781e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.806822233e-01 lpclm = -1.944471501e-7
+ pdiblc1 = 5.395309339e-01 lpdiblc1 = -2.029924265e-7
+ pdiblc2 = 1.009816291e-02 lpdiblc2 = -4.337771860e-9
+ pdiblcb = -7.427084443e-02 lpdiblcb = 2.516685754e-8
+ drout = -2.184018285e-01 ldrout = 6.223425964e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.757411360e-08 lalpha0 = 1.239108811e-15
+ alpha1 = 5.406994840e-01 lalpha1 = 1.579863734e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.422128596e-01 lkt1 = -1.458275149e-8
+ kt2 = -3.610075491e-02 lkt2 = -1.274268523e-10
+ at = 1.220672433e+05 lat = -3.674433855e-2
+ ute = -8.637901776e-01 lute = -1.849837664e-7
+ ua1 = 1.402279640e-09 lua1 = -1.576620366e-16
+ ub1 = -8.575982110e-19 lub1 = 9.084763742e-26
+ uc1 = -3.564555919e-12 luc1 = 2.184446813e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.60 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.262913778e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.765635388e-8
+ k1 = 2.050795932e-01 lk1 = 1.830701804e-7
+ k2 = 7.863177628e-02 lk2 = -5.890010271e-08 pk2 = 1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.618143394e-01 ldsub = 7.740536886e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446112e-03 lcdscd = -1.783892580e-09 wcdscd = 6.938893904e-24
+ cit = 0.0
+ voff = {-1.109742158e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.760456345e-8
+ nfactor = 4.519022990e+00 lnfactor = -7.883151319e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.525776721e-02 letab = -2.327665451e-08 wetab = -1.344410694e-23 petab = -1.951563910e-30
+ u0 = 2.458504396e-02 lu0 = -1.551688163e-9
+ ua = -1.881576616e-09 lua = 2.024024342e-16
+ ub = 2.589559975e-18 lub = -4.131032724e-25
+ uc = 6.187197712e-11 luc = 8.003006735e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.078372716e+04 lvsat = 2.929729196e-2
+ a0 = 1.5
+ ags = 9.337213088e-01 lags = 8.248105476e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.208158801e-02 lketa = -2.744240334e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.727091359e-01 lpclm = -1.392960087e-7
+ pdiblc1 = -8.200367215e-02 lpdiblc1 = 1.144787488e-7
+ pdiblc2 = -5.487871871e-03 lpdiblc2 = 3.623356504e-9
+ pdiblcb = 5.667376270e-02 lpdiblcb = -4.171781455e-08 ppdiblcb = 6.938893904e-30
+ drout = 1.518101815e+00 ldrout = -2.646391535e-7
+ pscbe1 = 8.089503007e+08 lpscbe1 = -4.571688292e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.876240960e-08 lalpha0 = -4.475716150e-15
+ alpha1 = 0.85
+ beta0 = 1.338015376e+01 lbeta0 = 2.450987415e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.018500067e-01 lkt1 = 1.587906831e-8
+ kt2 = -4.414385625e-02 lkt2 = 3.980876710e-9
+ at = 7.246399777e+04 lat = -1.140769520e-02 wat = -5.820766091e-17
+ ute = -1.128830784e+00 lute = -4.960473507e-8
+ ua1 = 2.259287292e-09 lua1 = -5.954095471e-16
+ ub1 = -2.127094562e-18 lub1 = 7.392886007e-25 wub1 = 7.703719778e-40
+ uc1 = -7.344148208e-11 luc1 = 5.753662374e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.61 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.364038796e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.029355277e-08 wvth0 = -4.358799651e-08 pvth0 = 1.136713926e-14
+ k1 = 0.90707349
+ k2 = -8.578994760e-02 lk2 = -1.602121903e-08 wk2 = -5.033029595e-08 pk2 = 1.312543656e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586434640e-01 ldsub = -3.511233284e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-9.930381000e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804189e-8
+ nfactor = -9.804248055e+00 lnfactor = 2.946993431e-06 wnfactor = 1.238450548e-05 pnfactor = -3.229705646e-12
+ eta0 = 6.941433251e-04 leta0 = -8.671466817e-16
+ etab = -0.043998
+ u0 = -4.408554454e-02 lu0 = 1.635663993e-08 wu0 = 3.886073989e-08 pu0 = -1.013433691e-14
+ ua = -7.946750893e-10 lua = -8.104626744e-17 wua = -3.912580058e-16 pua = 1.020346103e-22
+ ub = -5.749018091e-18 lub = 1.761481147e-24 wub = 5.122208891e-24 pub = -1.335800368e-30
+ uc = 3.967248006e-10 luc = -7.932192169e-17 wuc = -3.141523801e-16 puc = 8.192654260e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.010435078e+04 lvsat = 4.251376381e-02 wvsat = 8.676671606e-02 pvsat = -2.262754482e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.744150730e-01 lketa = 1.541941749e-07 wketa = 4.200474090e-07 pketa = -1.095424836e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.991951134e-01 lpclm = -4.188878082e-08 wpclm = 1.214906352e-07 ppclm = -3.168305679e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -7.983346087e-08 lalpha0 = 2.645242653e-14 walpha0 = 9.047174962e-14 palpha0 = -2.359376570e-20
+ alpha1 = 0.85
+ beta0 = 1.775146819e+01 lbeta0 = -8.948788635e-07 wbeta0 = -2.477202668e-06 pbeta0 = 6.460197750e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.824689802e-01 lkt1 = 6.298196792e-08 wkt1 = 2.154089277e-07 pkt1 = -5.617563261e-14
+ kt2 = -0.028878939
+ at = 1.830122700e+05 lat = -4.023713693e-02 wat = -2.154089277e-01 pat = 5.617563261e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.62 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.759269925e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.755409384e-09 wvth0 = -3.687103082e-08 pvth0 = 1.008563624e-14
+ k1 = 0.90707349
+ k2 = -2.991464838e-01 lk2 = 2.468422109e-08 wk2 = 1.675052933e-07 pk2 = -2.843454417e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.312030375e+01 lnfactor = -5.242410110e-06 wnfactor = -3.619665670e-05 pnfactor = 6.038899963e-12
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 7.925577053e-02 lu0 = -7.175156208e-09 wu0 = -5.758045052e-08 pu0 = 8.265292041e-15
+ ua = -1.940683164e-09 lua = 1.375960290e-16 wua = 9.743342244e-16 pua = -1.585012689e-22
+ ub = 3.831602461e-18 lub = -6.636712562e-26 wub = -2.280067920e-24 pub = 7.645041575e-32
+ uc = -5.553195725e-10 luc = 1.023148161e-16 wuc = 7.330222203e-16 puc = -1.178597107e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.614499104e+05 lvsat = 2.841298718e-04 wvsat = -3.011946282e-02 pvsat = -3.272982915e-10
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 8.508406928e-01 lketa = -1.368032716e-07 wketa = -9.801106209e-07 pketa = 1.575880663e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.796361268e-01 wpclm = -4.457530670e-8
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.132579954e-07 lalpha0 = -2.946532004e-14 walpha0 = -2.111007491e-13 palpha0 = 3.394204505e-20
+ alpha1 = 0.85
+ beta0 = 8.832221556e+00 lbeta0 = 8.067885250e-07 wbeta0 = 5.780139559e-06 pbeta0 = -9.293655192e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 2.153678204e-01 lkt1 = -7.015552391e-08 wkt1 = -5.026208312e-07 pkt1 = 8.081439297e-14
+ kt2 = -0.028878939
+ at = -3.956080734e+05 lat = 7.015552391e-02 wat = 5.026208312e-01 pat = -8.081439297e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.63 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.167023583e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.446859454e-06 wvth0 = 4.718153834e-08 pvth0 = -4.718662734e-12
+ k1 = 6.997665621e-01 lk1 = -1.317730536e-05 wk1 = -9.643851283e-08 pk1 = 9.644891469e-12
+ k2 = -7.901980754e-02 lk2 = 4.708863997e-06 wk2 = 3.446196536e-08 pk2 = -3.446568243e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.039000940e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.378218192e-07 wvoff = -3.204212391e-09 pvoff = 3.204557998e-13
+ nfactor = 4.940526918e+00 lnfactor = -1.018436755e-04 wnfactor = -7.453460580e-07 pnfactor = 7.454264510e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.405554935e-02 lu0 = 7.949608000e-07 wu0 = 5.817944959e-09 pu0 = -5.818572482e-13
+ ua = -1.591070566e-09 lua = 5.419837178e-14 wua = 3.966524436e-16 pua = -3.966952265e-20
+ ub = 1.361072919e-18 lub = -1.127350777e-23 wub = -8.250551188e-26 pub = 8.251441093e-30
+ uc = 8.024276129e-11 luc = -3.170918107e-15 wuc = -2.320646127e-17 puc = 2.320896432e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.353357948e+00 la0 = 9.243049175e-07 wa0 = 6.764553844e-09 pa0 = -6.765283469e-13
+ ags = 3.396356791e-01 lags = 5.244886534e-07 wags = 3.838486271e-09 pags = -3.838900291e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -3.424943097e-08 lb0 = 1.994758229e-12 wb0 = 1.459869918e-14 pb0 = -1.460027380e-18
+ b1 = 2.963064236e-08 lb1 = -1.725750355e-12 wb1 = -1.262995682e-14 pb1 = 1.263131909e-18
+ keta = -8.748251028e-03 lketa = 4.202104218e-07 wketa = 3.075322840e-09 pketa = -3.075654544e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.606981592e-02 lpclm = 9.295484095e-06 wpclm = 6.802928501e-08 ppclm = -6.803662265e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.093461422e-03 lpdiblc2 = 3.054118263e-07 wpdiblc2 = 2.235165804e-09 ppdiblc2 = -2.235406889e-13
+ pdiblcb = 3.033677576e+00 lpdiblcb = -3.059007485e-04 wpdiblcb = -2.238743995e-06 ppdiblcb = 2.238985466e-10
+ drout = 0.56
+ pscbe1 = -5.231123437e+08 lpscbe1 = 7.481930351e+04 wpscbe1 = 5.475673639e+02 ppscbe1 = -5.476264245e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.778741884e-01 lkt1 = -8.506729023e-07 wkt1 = -6.225675686e-09 pkt1 = 6.226347188e-13
+ kt2 = -4.190194228e-02 lkt2 = 1.238534702e-06 wkt2 = 9.064254145e-09 pkt2 = -9.065231815e-13
+ at = 2.238038370e+05 lat = -4.880910095e+00 wat = -3.572109000e-02 pat = 3.572494288e-6
+ ute = -8.751456826e-01 lute = -2.402802313e-05 wute = -1.758498231e-07 pute = 1.758687902e-11
+ ua1 = 7.966636434e-10 lua1 = 3.243713395e-14 wua1 = 2.373921581e-16 pua1 = -2.374177633e-20
+ ub1 = -4.993223950e-20 lub1 = -5.195937978e-23 wub1 = -3.802663121e-25 pub1 = 3.803073276e-29
+ uc1 = 1.150093803e-10 luc1 = -8.119977561e-15 wuc1 = -5.942630444e-17 puc1 = 5.943271416e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.64 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {8.800473258e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.825037535e-06 wvth0 = -3.145435889e-07 pvth0 = 2.519741379e-12
+ k1 = -2.473051351e-01 lk1 = 5.774343698e-06 wk1 = 6.429234189e-07 pk1 = -5.150321923e-12
+ k2 = 2.594129521e-01 lk2 = -2.063441530e-06 wk2 = -2.297464358e-07 pk2 = 1.840449531e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.353669715e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.918551322e-07 wvoff = 2.136141594e-08 pvoff = -1.711217318e-13
+ nfactor = -2.379123037e+00 lnfactor = 4.462827335e-05 wnfactor = 4.968973720e-06 pnfactor = -3.980538511e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 7.119051385e-02 lu0 = -3.483547477e-07 wu0 = -3.878629973e-08 pu0 = 3.107087468e-13
+ ua = 2.304243578e-09 lua = -2.374992594e-14 wua = -2.644349624e-15 pua = 2.118331895e-20
+ ub = 5.508298653e-19 lub = 4.940092589e-24 wub = 5.500367459e-25 pub = -4.406226663e-30
+ uc = -1.476556376e-10 luc = 1.389507982e-15 wuc = 1.547097418e-16 puc = -1.239346634e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.419789058e+00 la0 = -4.050338160e-07 wa0 = -4.509702563e-08 pa0 = 3.612626215e-13
+ ags = 3.773314254e-01 lags = -2.298328578e-07 wags = -2.558990848e-08 pags = 2.049952806e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.091166829e-07 lb0 = -8.741103958e-13 wb0 = -9.732466122e-14 pb0 = 7.796470336e-19
+ b1 = -9.440149266e-08 lb1 = 7.562301558e-13 wb1 = 8.419971215e-14 pb1 = -6.745058753e-19
+ keta = 2.145287025e-02 lketa = -1.841377530e-07 wketa = -2.050215227e-08 pketa = 1.642383543e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.920098602e-01 lpclm = -4.073315334e-06 wpclm = -4.535285667e-07 ppclm = 3.633120293e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.985692136e-02 lpdiblc2 = -1.338325861e-07 wpdiblc2 = -1.490110536e-08 ppdiblc2 = 1.193695662e-13
+ pdiblcb = -1.895184474e+01 lpdiblcb = 1.340468336e-04 wpdiblcb = 1.492495997e-05 ppdiblcb = -1.195606604e-10
+ drout = 0.56
+ pscbe1 = 4.854257521e+09 lpscbe1 = -3.278609410e+04 wpscbe1 = -3.650449093e+03 ppscbe1 = 2.924296649e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.390132610e-01 lkt1 = 3.727679960e-07 wkt1 = 4.150450457e-08 pkt1 = -3.324837042e-13
+ kt2 = 4.711331008e-02 lkt2 = -5.427304638e-07 wkt2 = -6.042836096e-08 pkt2 = 4.840786680e-13
+ at = -1.269941207e+05 lat = 2.138832764e+00 wat = 2.381406000e-01 pat = -1.907693385e-6
+ ute = -2.602073914e+00 lute = 1.052916815e-05 wute = 1.172332154e-06 pute = -9.391302005e-12
+ ua1 = 3.127966642e-09 lua1 = -1.421407145e-14 wua1 = -1.582614388e-15 pua1 = 1.267798518e-20
+ ub1 = -3.784326840e-18 lub1 = 2.276879141e-23 wub1 = 2.535108747e-24 pub1 = -2.030821366e-29
+ uc1 = -4.685849676e-10 luc1 = 3.558204046e-15 wuc1 = 3.961753629e-16 puc1 = -3.173676051e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.65 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.170743503e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.266129549e-8
+ k1 = 4.567336080e-01 lk1 = 1.344399904e-7
+ k2 = 1.114140034e-02 lk2 = -7.459125980e-08 wk2 = -1.734723476e-24 pk2 = -2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.168391204e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.343248247e-8
+ nfactor = 3.469646930e+00 lnfactor = -2.224971222e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.811640691e-02 lu0 = -3.297294898e-9
+ ua = -6.221534367e-10 lua = -3.071857119e-16
+ ub = 1.157713655e-18 lub = 7.847642182e-26
+ uc = 2.622213792e-11 luc = -3.389667350e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.501305188e+00 la0 = -1.058042092e-6
+ ags = 3.581621046e-01 lags = -7.627153156e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.285724033e-02 lketa = 9.071320047e-08 wketa = -1.734723476e-24 pketa = -2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.673104246e-01 lpclm = 3.611594172e-06 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.955579854e-03 lpdiblc2 = 1.560443807e-9
+ pdiblcb = -4.418017311e+00 lpdiblcb = 1.761945233e-5
+ drout = 0.56
+ pscbe1 = 7.778430133e+08 lpscbe1 = -1.308098334e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912466833e-01 lkt1 = -9.879836114e-9
+ kt2 = -2.057476356e-02 lkt2 = -4.957910604e-10
+ at = 140000.0
+ ute = -1.490445232e+00 lute = 1.624148668e-6
+ ua1 = 1.251425227e-09 lua1 = 8.185002439e-16
+ ub1 = -9.358332547e-19 lub1 = -4.988112379e-26
+ uc1 = -3.054834705e-11 luc1 = 4.918641870e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.66 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.106045433e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.086103068e-7
+ k1 = 4.408190516e-01 lk1 = 1.982698706e-7
+ k2 = 1.863132370e-02 lk2 = -1.046317395e-07 wk2 = 6.938893904e-24 pk2 = -1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.606520361e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.999511228e-8
+ nfactor = 3.549780143e+00 lnfactor = -2.546368387e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.933554941e-02 lu0 = -8.187014548e-9
+ ua = -2.414911465e-10 lua = -1.833940696e-15
+ ub = 6.589395849e-19 lub = 2.078952480e-24
+ uc = -3.494870781e-12 luc = 1.157988951e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.515523305e+00 la0 = -1.115067914e-6
+ ags = 1.366518094e-01 lags = 8.121588595e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.846356849e-02 lketa = -7.501572108e-08 pketa = -2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.091009455e-01 lpclm = 9.649571892e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.381838483e-03 lpdiblc2 = 7.872383663e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.901616173e+08 lpscbe1 = 2.208614822e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.957509478e-01 lkt1 = 8.185804823e-9
+ kt2 = -2.371415082e-02 lkt2 = 1.209561941e-8
+ at = 1.689553184e+05 lat = -1.161335857e-1
+ ute = -1.752105721e+00 lute = 2.673612892e-6
+ ua1 = -7.113229936e-10 lua1 = 8.690663327e-15
+ ub1 = 8.493023065e-19 lub1 = -7.209677841e-24
+ uc1 = -6.285819551e-12 luc1 = -4.812538692e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.67 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.342275017e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.110959292e-8
+ k1 = 6.002258295e-01 lk1 = -1.222630466e-7
+ k2 = -5.139249434e-02 lk2 = 3.617117345e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.000814656e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.181140900e-8
+ nfactor = 2.759531280e+00 lnfactor = -9.573470380e-7
+ eta0 = 1.583042774e-01 leta0 = -1.574531447e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 2.787667965e-02 lu0 = -5.253539668e-9
+ ua = -9.177990006e-10 lua = -4.740303314e-16
+ ub = 1.500559190e-18 lub = 3.866355608e-25
+ uc = 3.787088470e-11 luc = 3.262121312e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.989214000e+04 lvsat = 2.032474338e-2
+ a0 = 1.430132279e+00 la0 = -9.433648340e-7
+ ags = 3.661307571e-01 lags = 3.507258042e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.742407017e-02 lketa = 3.736236032e-08 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.244546611e-01 lpclm = 2.667012826e-7
+ pdiblc1 = 4.418486520e-01 lpdiblc1 = -1.042565435e-7
+ pdiblc2 = 4.781655300e-03 lpdiblc2 = 1.036079606e-9
+ pdiblcb = -3.645777836e-04 lpdiblcb = -4.953656210e-8
+ drout = 7.244550742e-01 ldrout = -3.306839609e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.121294320e-08 lalpha0 = -2.438969205e-15
+ alpha1 = 1.004650258e+00 lalpha1 = -3.109685737e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.270979414e-01 lkt1 = 7.121790080e-8
+ kt2 = 1.029101439e-03 lkt2 = -3.765776583e-8
+ at = 1.369598812e+05 lat = -5.179760850e-02 wat = -1.164153218e-16
+ ute = 2.085940234e-01 lute = -1.268934703e-6
+ ua1 = 6.000602418e-09 lua1 = -4.805582324e-15
+ ub1 = -4.725912025e-18 lub1 = 4.000885084e-24 pub1 = 3.081487911e-45
+ uc1 = -7.900628978e-11 luc1 = 9.809991654e-17 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.68 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.977095171e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.057139584e-9
+ k1 = 3.932297063e-01 lk1 = 8.696573668e-8
+ k2 = 5.920903785e-03 lk2 = -2.176040699e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.054929839e-01 ldsub = 5.509492874e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.573674280e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.092439875e-9
+ nfactor = 6.240200030e-01 lnfactor = 1.201197864e-6
+ eta0 = -4.954530748e-01 leta0 = 5.033556343e-07 weta0 = -1.040834086e-22 peta0 = 1.127570259e-28
+ etab = -1.702508962e-01 letab = 8.680215367e-8
+ u0 = 2.383561950e-02 lu0 = -1.168892645e-9
+ ua = -1.286096305e-09 lua = -1.017605720e-16
+ ub = 1.987544147e-18 lub = -1.056020158e-25
+ uc = 6.258845349e-11 luc = 7.637040637e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.060478235e+04 lvsat = 6.003585447e-2
+ a0 = -5.279722970e-01 la0 = 1.035859858e-6
+ ags = 3.227856408e-01 lags = 3.945384409e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.161186290e-02 lketa = -4.252605433e-08 wketa = -1.387778781e-23 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.806822233e-01 lpclm = -1.944471501e-7
+ pdiblc1 = 5.395309339e-01 lpdiblc1 = -2.029924265e-7
+ pdiblc2 = 1.009816291e-02 lpdiblc2 = -4.337771860e-9
+ pdiblcb = -7.427084443e-02 lpdiblcb = 2.516685754e-8
+ drout = -2.184018285e-01 ldrout = 6.223425964e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.757411360e-08 lalpha0 = 1.239108811e-15
+ alpha1 = 5.406994840e-01 lalpha1 = 1.579863734e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.422128596e-01 lkt1 = -1.458275149e-8
+ kt2 = -3.610075491e-02 lkt2 = -1.274268523e-10
+ at = 1.220672433e+05 lat = -3.674433855e-2
+ ute = -8.637901776e-01 lute = -1.849837664e-7
+ ua1 = 1.402279640e-09 lua1 = -1.576620366e-16
+ ub1 = -8.575982110e-19 lub1 = 9.084763742e-26
+ uc1 = -3.564555919e-12 luc1 = 2.184446813e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.69 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.262913778e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.765635388e-8
+ k1 = 2.050795932e-01 lk1 = 1.830701804e-7
+ k2 = 7.863177628e-02 lk2 = -5.890010271e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.618143394e-01 ldsub = 7.740536886e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446112e-03 lcdscd = -1.783892580e-09 wcdscd = 6.938893904e-24
+ cit = 0.0
+ voff = {-1.109742158e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.760456345e-8
+ nfactor = 4.519022990e+00 lnfactor = -7.883151319e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.525776721e-02 letab = -2.327665451e-08 wetab = 4.336808690e-25 petab = -4.770489559e-30
+ u0 = 2.458504396e-02 lu0 = -1.551688163e-9
+ ua = -1.881576616e-09 lua = 2.024024342e-16
+ ub = 2.589559975e-18 lub = -4.131032724e-25
+ uc = 6.187197712e-11 luc = 8.003006735e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.078372716e+04 lvsat = 2.929729196e-2
+ a0 = 1.5
+ ags = 9.337213088e-01 lags = 8.248105476e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.208158801e-02 lketa = -2.744240334e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.727091359e-01 lpclm = -1.392960087e-7
+ pdiblc1 = -8.200367215e-02 lpdiblc1 = 1.144787488e-7
+ pdiblc2 = -5.487871871e-03 lpdiblc2 = 3.623356504e-09 wpdiblc2 = 1.734723476e-24 ppdiblc2 = 8.673617380e-31
+ pdiblcb = 5.667376270e-02 lpdiblcb = -4.171781455e-08 ppdiblcb = 6.938893904e-30
+ drout = 1.518101815e+00 ldrout = -2.646391535e-7
+ pscbe1 = 8.089503007e+08 lpscbe1 = -4.571688292e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.876240960e-08 lalpha0 = -4.475716150e-15
+ alpha1 = 0.85
+ beta0 = 1.338015376e+01 lbeta0 = 2.450987415e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.018500067e-01 lkt1 = 1.587906831e-8
+ kt2 = -4.414385625e-02 lkt2 = 3.980876710e-9
+ at = 7.246399777e+04 lat = -1.140769520e-2
+ ute = -1.128830784e+00 lute = -4.960473507e-8
+ ua1 = 2.259287292e-09 lua1 = -5.954095471e-16
+ ub1 = -2.127094562e-18 lub1 = 7.392886007e-25 pub1 = 1.925929944e-46
+ uc1 = -7.344148208e-11 luc1 = 5.753662374e-17 puc1 = 1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.70 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.875346872e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.549151562e-9
+ k1 = 0.90707349
+ k2 = -1.422183479e-01 lk2 = -1.305482221e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586434640e-01 ldsub = -3.511233285e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-9.930381000e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804189e-8
+ nfactor = 4.080785197e+00 lnfactor = -6.740288509e-7
+ eta0 = 6.941433251e-04 leta0 = -8.671466817e-16
+ etab = -0.043998
+ u0 = -5.163712314e-04 lu0 = 4.994409498e-9
+ ua = -1.233338581e-09 lua = 3.335102999e-17
+ ub = -6.193647714e-21 lub = 2.638329318e-25
+ uc = 4.450918314e-11 luc = 1.253098032e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.373838699e+05 lvsat = 1.714462714e-2
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.034740047e-01 lketa = 3.137933746e-08 pketa = 2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.354057609e-01 lpclm = -7.741061073e-8
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.16e-8
+ alpha1 = 0.85
+ beta0 = 1.497412343e+01 lbeta0 = -1.705862324e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.24096074
+ kt2 = -0.028878939
+ at = -5.849597014e+04 lat = 2.274483099e-2
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.71 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {7.299937748e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.472835104e-08 wvth0 = -1.742881241e-07 pvth0 = 3.325173404e-14
+ k1 = 0.90707349
+ k2 = 1.769009749e-02 lk2 = -3.181377489e-08 wk2 = -1.150913923e-07 pk2 = 2.195782638e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587461769e-01 ldsub = -2.310740521e-11 wdsub = -1.080280217e-10 pdsub = 2.061023415e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = -6.481886456e+00 lnfactor = 1.341181023e-06 wnfactor = -8.741959909e-07 pnfactor = 1.667843563e-13
+ eta0 = -1.632446765e-02 leta0 = 3.246912159e-09 weta0 = 1.517944113e-08 peta0 = -2.896024855e-15
+ etab = -0.043998
+ u0 = 3.603765658e-02 lu0 = -1.979587253e-09 wu0 = -1.903283172e-08 pu0 = 3.631197832e-15
+ ua = -2.620746877e-09 lua = 2.980491091e-16 wua = 1.580904812e-15 pua = -3.016145055e-22
+ ub = 1.618074477e-17 lub = -2.824408301e-24 wub = -1.329466311e-23 pub = 2.536435597e-30
+ uc = 1.680052029e-10 luc = -1.103033130e-17 wuc = 8.786570671e-17 puc = -1.676354672e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.896559766e+05 lvsat = -1.263783590e-01 wvsat = -5.904365558e-01 pvsat = 1.126470287e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.635612593e-06 lb0 = 1.075195984e-12 wb0 = 5.026583212e-12 pb0 = -9.590017046e-19
+ b1 = 3.860048929e-06 lb1 = -7.364432949e-13 wb1 = -3.442901161e-12 pb1 = 6.568573409e-19
+ keta = -9.099966544e-01 lketa = 1.661739677e-07 wketa = 5.904365558e-07 pketa = -1.126470287e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 9.092221223e-02 lpclm = 7.390627578e-09 wpclm = 3.455147252e-08 ppclm = -6.591937237e-15
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.342008000e-08 lalpha0 = 8.589200983e-15
+ alpha1 = 0.85
+ beta0 = 2.021621011e+01 lbeta0 = -1.170702981e-06 wbeta0 = -4.373604117e-06 pbeta0 = 8.344224351e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.385031506e-01 lkt1 = 1.140027264e-07 wkt1 = 4.373604117e-07 pkt1 = -8.344224351e-14
+ kt2 = -0.028878939
+ at = 4.866397872e+05 lat = -8.125943962e-02 wat = -2.842842676e-01 pat = 5.423745828e-8
+ ute = -9.316384008e-02 lute = -2.338806196e-07 wute = -1.093401029e-06 pute = 2.086056088e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.72 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.73 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.503030477e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.175519114e-7
+ k1 = 6.310871457e-01 lk1 = -1.262268888e-6
+ k2 = -5.447745820e-02 lk2 = 4.510673736e-07 wk2 = -2.775557562e-23 pk2 = 2.220446049e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.061819981e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.193944404e-8
+ nfactor = 4.409723085e+00 lnfactor = -9.755720117e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.819884287e-02 lu0 = 7.615018832e-8
+ ua = -1.308591527e-09 lua = 5.191722935e-15
+ ub = 1.302315995e-18 lub = -1.079901978e-24
+ uc = 6.371610434e-11 luc = -3.037458086e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.358175376e+00 la0 = 8.854020668e-8
+ ags = 3.423692862e-01 lags = 5.024135747e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.385285691e-08 lb0 = 1.910801322e-13
+ b1 = 2.063612306e-08 lb1 = -1.653115657e-13
+ keta = -6.558136603e-03 lketa = 4.025242849e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.762224597e-02 lpclm = 8.904248667e-07 ppclm = 2.220446049e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -5.016711857e-04 lpdiblc2 = 2.925574203e-08 ppdiblc2 = -1.387778781e-29
+ pdiblcb = 1.439339104e+00 lpdiblcb = -2.930257643e-05 wpdiblcb = -2.498001805e-22 ppdiblcb = -5.329070518e-27
+ drout = 0.56
+ pscbe1 = -1.331581032e+08 lpscbe1 = 7.167025156e+03 ppscbe1 = 1.907348633e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.823078504e-01 lkt1 = -8.148691321e-8
+ kt2 = -3.544676512e-02 lkt2 = 1.186406308e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.000378464e+00 lute = -2.301671335e-6
+ ua1 = 9.657242647e-10 lua1 = 3.107189510e-15
+ ub1 = -3.207417704e-19 lub1 = -4.977247376e-24
+ uc1 = 7.268848809e-11 luc1 = -7.778217749e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.74 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.170743503e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.266129549e-8
+ k1 = 4.567336080e-01 lk1 = 1.344399904e-7
+ k2 = 1.114140034e-02 lk2 = -7.459125980e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.168391204e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.343248247e-8
+ nfactor = 3.469646930e+00 lnfactor = -2.224971222e-06 wnfactor = -3.552713679e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.811640691e-02 lu0 = -3.297294898e-9
+ ua = -6.221534367e-10 lua = -3.071857119e-16
+ ub = 1.157713655e-18 lub = 7.847642182e-26
+ uc = 2.622213792e-11 luc = -3.389667350e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.501305188e+00 la0 = -1.058042092e-6
+ ags = 3.581621046e-01 lags = -7.627153156e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.285724033e-02 lketa = 9.071320047e-08 wketa = -3.469446952e-24
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.673104246e-01 lpclm = 3.611594172e-06 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.955579854e-03 lpdiblc2 = 1.560443807e-9
+ pdiblcb = -4.418017311e+00 lpdiblcb = 1.761945233e-5
+ drout = 0.56
+ pscbe1 = 7.778430133e+08 lpscbe1 = -1.308098334e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912466833e-01 lkt1 = -9.879836114e-9
+ kt2 = -2.057476356e-02 lkt2 = -4.957910604e-10
+ at = 140000.0
+ ute = -1.490445232e+00 lute = 1.624148668e-6
+ ua1 = 1.251425227e-09 lua1 = 8.185002439e-16
+ ub1 = -9.358332547e-19 lub1 = -4.988112379e-26
+ uc1 = -3.054834705e-11 luc1 = 4.918641870e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.75 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.106045433e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.086103068e-7
+ k1 = 4.408190516e-01 lk1 = 1.982698706e-7
+ k2 = 1.863132370e-02 lk2 = -1.046317395e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.606520361e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.999511228e-8
+ nfactor = 3.549780143e+00 lnfactor = -2.546368387e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.933554941e-02 lu0 = -8.187014548e-9
+ ua = -2.414911465e-10 lua = -1.833940696e-15
+ ub = 6.589395849e-19 lub = 2.078952480e-24
+ uc = -3.494870781e-12 luc = 1.157988951e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.515523305e+00 la0 = -1.115067914e-6
+ ags = 1.366518094e-01 lags = 8.121588595e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.846356849e-02 lketa = -7.501572108e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.091009455e-01 lpclm = 9.649571892e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.381838483e-03 lpdiblc2 = 7.872383663e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.901616173e+08 lpscbe1 = 2.208614822e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.957509478e-01 lkt1 = 8.185804823e-9
+ kt2 = -2.371415082e-02 lkt2 = 1.209561941e-8
+ at = 1.689553184e+05 lat = -1.161335857e-1
+ ute = -1.752105721e+00 lute = 2.673612892e-6
+ ua1 = -7.113229936e-10 lua1 = 8.690663327e-15
+ ub1 = 8.493023065e-19 lub1 = -7.209677841e-24 pub1 = -3.081487911e-45
+ uc1 = -6.285819551e-12 luc1 = -4.812538692e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.76 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.342275017e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.110959292e-8
+ k1 = 6.002258295e-01 lk1 = -1.222630466e-7
+ k2 = -5.139249434e-02 lk2 = 3.617117345e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.000814656e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.181140900e-8
+ nfactor = 2.759531280e+00 lnfactor = -9.573470380e-7
+ eta0 = 1.583042774e-01 leta0 = -1.574531447e-7
+ etab = -5.546995125e-02 letab = -2.921681861e-8
+ u0 = 2.787667965e-02 lu0 = -5.253539668e-9
+ ua = -9.177990006e-10 lua = -4.740303314e-16
+ ub = 1.500559190e-18 lub = 3.866355608e-25
+ uc = 3.787088470e-11 luc = 3.262121312e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.989214000e+04 lvsat = 2.032474338e-2
+ a0 = 1.430132279e+00 la0 = -9.433648340e-7
+ ags = 3.661307571e-01 lags = 3.507258042e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.742407017e-02 lketa = 3.736236032e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.244546611e-01 lpclm = 2.667012826e-7
+ pdiblc1 = 4.418486520e-01 lpdiblc1 = -1.042565435e-07 wpdiblc1 = 4.440892099e-22
+ pdiblc2 = 4.781655300e-03 lpdiblc2 = 1.036079606e-9
+ pdiblcb = -3.645777836e-04 lpdiblcb = -4.953656210e-8
+ drout = 7.244550742e-01 ldrout = -3.306839609e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.121294320e-08 lalpha0 = -2.438969205e-15
+ alpha1 = 1.004650258e+00 lalpha1 = -3.109685737e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.270979414e-01 lkt1 = 7.121790080e-8
+ kt2 = 1.029101439e-03 lkt2 = -3.765776583e-8
+ at = 1.369598812e+05 lat = -5.179760850e-02 wat = 1.164153218e-16
+ ute = 2.085940234e-01 lute = -1.268934703e-6
+ ua1 = 6.000602418e-09 lua1 = -4.805582324e-15
+ ub1 = -4.725912025e-18 lub1 = 4.000885084e-24 pub1 = -3.081487911e-45
+ uc1 = -7.900628978e-11 luc1 = 9.809991654e-17 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.77 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.236711974e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.929884253e-08 wvth0 = -1.900218456e-08 pvth0 = 1.920714212e-14
+ k1 = -1.781222905e-01 lk1 = 6.644803362e-07 wk1 = 4.181908098e-07 pk1 = -4.227014158e-13
+ k2 = 1.938136854e-01 lk2 = -2.116798002e-07 wk2 = -1.375247395e-07 pk2 = 1.390080813e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.858104465e-01 ldsub = 7.498976201e-08 wdsub = 1.440627898e-08 pdsub = -1.456166511e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.457251973e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.675363950e-09 wvoff = -8.521321219e-09 pvoff = 8.613232189e-15
+ nfactor = -4.413252793e-01 lnfactor = 2.278033960e-06 wnfactor = 7.797603032e-07 pnfactor = -7.881707978e-13
+ eta0 = -4.954530747e-01 leta0 = 5.033556341e-07 weta0 = -9.483244051e-17 peta0 = 9.585536531e-23
+ etab = -1.722682838e-01 letab = 8.884130080e-08 wetab = 1.476590533e-09 petab = -1.492517039e-15
+ u0 = 4.889606133e-03 lu0 = 1.798147243e-08 wu0 = 1.386719346e-08 pu0 = -1.401676501e-14
+ ua = -1.982656674e-09 lua = 6.023128972e-16 wua = 5.098348240e-16 pua = -5.153339024e-22
+ ub = 1.028495504e-18 lub = 8.637909260e-25 wub = 7.019583914e-25 pub = -7.095297147e-31
+ uc = -9.882192274e-11 luc = 1.707883892e-16 wuc = 1.181414195e-16 puc = -1.194156928e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.562863936e+06 lvsat = -1.488750246e+00 wvsat = -1.121509507e+00 pvsat = 1.133606108e-6
+ a0 = -1.272953194e+00 la0 = 1.788876119e-06 wa0 = 5.452753582e-07 pa0 = -5.511566982e-13
+ ags = -5.738737879e+00 lags = 6.521441554e-06 wags = 4.436623033e-06 pags = -4.484476449e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.480044889e-17 lb0 = 1.496008653e-23 wb0 = 1.083292215e-23 pb0 = -1.094976605e-29
+ b1 = -8.560766018e-17 lb1 = 8.653102440e-23 wb1 = 6.265898593e-23 pb1 = -6.333482575e-29
+ keta = 2.099747374e-01 lketa = -2.025970308e-07 wketa = -1.159108555e-07 pketa = 1.171610700e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.695849122e-01 lpclm = 1.200056566e-07 wpclm = 2.277020771e-07 ppclm = -2.301580717e-13
+ pdiblc1 = -1.646971660e-01 lpdiblc1 = 5.088314777e-07 wpdiblc1 = 5.154470816e-07 ppdiblc1 = -5.210066939e-13
+ pdiblc2 = 3.137653477e-05 lpdiblc2 = 5.837594878e-09 wpdiblc2 = 7.368203088e-09 ppdiblc2 = -7.447676527e-15
+ pdiblcb = -5.236170481e-01 lpdiblcb = 4.793597093e-07 wpdiblcb = 3.288908655e-07 ppdiblcb = -3.324382824e-13
+ drout = -2.184024743e-01 ldrout = 6.223432491e-07 wdrout = 4.726609921e-13 pdrout = -4.777591138e-19
+ pscbe1 = -1.543739537e+09 lpscbe1 = 2.369019111e+03 wpscbe1 = 1.715457967e+03 ppscbe1 = -1.733960896e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.501090235e-05 lalpha0 = -2.525155931e-11 walpha0 = -1.828609740e-11 palpha0 = 1.848333125e-17
+ alpha1 = 5.406994840e-01 lalpha1 = 1.579863734e-7
+ beta0 = 4.070255265e+01 lbeta0 = -2.713207642e-05 wbeta0 = -1.964692325e-05 pbeta0 = 1.985883496e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.950657684e-01 lkt1 = 3.884022869e-08 wkt1 = 3.868473517e-08 pkt1 = -3.910198873e-14
+ kt2 = -3.847883851e-02 lkt2 = 2.276306765e-09 wkt2 = 1.740595491e-09 pkt2 = -1.759369554e-15
+ at = -1.327699865e+05 lat = 2.208415655e-01 wat = 1.865235232e-01 pat = -1.885353659e-7
+ ute = -1.408217571e+00 lute = 3.653158208e-07 wute = 3.984838308e-07 pute = -4.027818774e-13
+ ua1 = -2.887400415e-10 lua1 = 1.551596983e-15 wua1 = 1.237711418e-15 pua1 = -1.251061373e-21
+ ub1 = -5.486267437e-19 lub1 = -2.214563962e-25 wub1 = -2.261461040e-25 pub1 = 2.285853159e-31
+ uc1 = -2.195792942e-10 luc1 = 2.401891414e-16 wuc1 = 1.581080994e-16 puc1 = -1.598134534e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.78 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.551590434e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.696206559e-09 wvth0 = 5.206403179e-08 pvth0 = -1.709248626e-14
+ k1 = 1.347783586e+00 lk1 = -1.149310229e-07 wk1 = -8.363816188e-07 pk1 = 2.181166167e-13
+ k2 = -2.966823963e-01 lk2 = 3.885873141e-08 wk2 = 2.747044530e-07 pk2 = -7.155281897e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.011794144e-01 ldsub = 6.713950838e-08 wdsub = -2.881255807e-08 pdsub = 7.513911793e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446104e-03 lcdscd = -1.783892576e-09 wcdscd = 5.922227986e-18 pcdscd = -3.024993450e-24
+ cit = 0.0
+ voff = {-1.342586770e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.153230201e-08 wvoff = 1.704264226e-08 pvoff = -4.444482458e-15
+ nfactor = 6.649713556e+00 lnfactor = -1.343969402e-06 wnfactor = -1.559520608e-06 pnfactor = 4.067011416e-13
+ eta0 = 1.000416472e+00 leta0 = -2.607135882e-07 weta0 = -7.090861232e-17 peta0 = 8.363554294e-23
+ etab = 4.929254235e-02 letab = -2.432886737e-08 wetab = -2.953181039e-09 petab = 7.701482633e-16
+ u0 = 7.336237544e-02 lu0 = -1.699345951e-08 wu0 = -3.570168978e-08 pu0 = 1.130232659e-14
+ ua = -4.884558750e-10 lua = -1.609039523e-16 wua = -1.019669650e-15 pua = 2.659155701e-22
+ ub = 4.507657262e-18 lub = -9.133161921e-25 wub = -1.403916784e-24 pub = 3.661218427e-31
+ uc = 3.846927297e-10 luc = -7.618412607e-17 wuc = -2.362828391e-16 puc = 6.161925649e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.515487836e+06 lvsat = 5.944147421e-01 wvsat = 1.907613558e+00 pvsat = -4.136275455e-7
+ a0 = 2.989961792e+00 la0 = -3.885611752e-07 wa0 = -1.090550714e-06 pa0 = 2.844003581e-13
+ ags = 1.305676835e+01 lags = -3.079039890e-06 wags = -8.873246066e-06 pags = 2.314018348e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.960089777e-17 lb0 = -7.719499726e-24 wb0 = -2.166584431e-23 pb0 = 5.650148874e-30
+ b1 = 1.712153204e-16 lb1 = -4.465055854e-23 wb1 = -1.253179719e-22 pb1 = 3.268117261e-29
+ keta = -2.946441610e-01 lketa = 5.515523782e-08 wketa = 2.318217109e-07 pketa = -6.045585669e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.394903759e+00 lpclm = -3.015556556e-07 wpclm = -4.554041545e-07 ppclm = 1.187630279e-13
+ pdiblc1 = 1.326452528e+00 lpdiblc1 = -2.528269100e-07 wpdiblc1 = -1.030894164e-06 ppdiblc1 = 2.688427654e-13
+ pdiblc2 = 1.464570088e-02 lpdiblc2 = -1.627197395e-09 wpdiblc2 = -1.473640617e-08 ppdiblc2 = 3.843048417e-15
+ pdiblcb = 9.553661700e-01 lpdiblcb = -2.760842127e-07 wpdiblcb = -6.577817310e-07 ppdiblcb = 1.715402665e-13
+ drout = 1.518103104e+00 ldrout = -2.646394890e-07 wdrout = -9.435148982e-13 pdrout = 2.456037045e-19
+ pscbe1 = 5.496429374e+09 lpscbe1 = -1.227000606e+03 wpscbe1 = -3.430915933e+03 ppscbe1 = 8.947348424e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -4.992789407e-05 lalpha0 = 1.302612876e-11 walpha0 = 3.657219481e-11 palpha0 = -9.537516395e-18
+ alpha1 = 0.85
+ beta0 = -4.030495154e+01 lbeta0 = 1.424542261e-05 wbeta0 = 3.929384649e-05 pbeta0 = -1.024728505e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.961441894e-01 lkt1 = -1.168752896e-08 wkt1 = -7.736947029e-08 pkt1 = 2.017687467e-14
+ kt2 = -3.938768905e-02 lkt2 = 2.740534894e-09 wkt2 = -3.481190971e-09 pkt2 = 9.078458658e-16
+ at = 5.821384572e+05 lat = -1.443236588e-01 wat = -3.730470465e-01 pat = 9.728544706e-8
+ ute = -3.997599746e-02 lute = -3.335628195e-07 wute = -7.969676618e-07 pute = 2.078380087e-13
+ ua1 = 5.641326653e-09 lua1 = -1.477398063e-15 wua1 = -2.475422833e-15 pua1 = 6.455556185e-22
+ ub1 = -2.745037501e-18 lub1 = 9.004394689e-25 wub1 = 4.522922110e-25 pub1 = -1.179514773e-31
+ uc1 = 3.585879945e-10 luc1 = -5.513061536e-17 wuc1 = -3.162161989e-16 puc1 = 8.246475765e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.79 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {1.197330485e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.617731150e-07 wvth0 = -4.463290577e-07 pvth0 = 1.128814540e-13
+ k1 = 9.070734932e-01 lk1 = -6.073390679e-16 wk1 = -2.329997528e-15 pk1 = 4.445310786e-22
+ k2 = -6.408110130e-02 lk2 = -2.180042990e-08 wk2 = -5.719115118e-08 pk2 = 1.500090805e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587285471e-01 ldsub = -2.569974795e-11 wdsub = -6.227504236e-11 pdsub = 1.624048392e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000032e-03 lcdscd = -6.426701185e-18 wcdscd = -2.371471769e-17 pcdscd = 4.703908270e-24
+ cit = 0.0
+ voff = {-9.930381134e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804160e-08 wvoff = 9.804734802e-16 pvoff = -2.105716712e-22
+ nfactor = 2.776520619e+01 lnfactor = -6.850594264e-06 wnfactor = -1.733538563e-05 pnfactor = 4.520825876e-12
+ eta0 = -1.126128123e-02 leta0 = 3.117806392e-09 weta0 = 8.750557806e-09 peta0 = -2.282022903e-15
+ etab = -4.399799986e-02 letab = -2.622341233e-17 wetab = -1.006036365e-16 petab = 1.919375769e-23
+ u0 = -3.519381827e-02 lu0 = 1.131647602e-08 wu0 = 2.538153316e-08 pu0 = -4.627322791e-15
+ ua = -1.822370922e-09 lua = 1.869624172e-16 wua = 4.311316193e-16 pua = -1.124330899e-22
+ ub = 8.025675296e-19 lub = 5.291933898e-26 wub = -5.919581861e-25 pub = 1.543744078e-31
+ uc = -5.270664684e-10 luc = 1.615899082e-16 wuc = 4.183545098e-16 puc = -1.091009992e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.200529879e+05 lvsat = 4.795466975e-02 wvsat = 4.080058742e-01 pvsat = -2.255085611e-8
+ a0 = 1.500000010e+00 la0 = -1.855308795e-15 wa0 = -7.117712642e-15 pa0 = 1.357959967e-21
+ ags = 1.250000002e+00 lags = -3.972386864e-16 wags = -1.523968507e-15 pags = 2.907523111e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.673484566e-07 lb0 = 6.972073460e-14 wb0 = 1.956808905e-13 pb0 = -5.103083672e-20
+ b1 = 1.831174339e-07 lb1 = -4.775446311e-14 wb1 = -1.340295096e-13 pb1 = 3.495301970e-20
+ keta = 3.206758066e-03 lketa = -2.252011195e-08 wketa = -1.512762640e-07 pketa = 3.945073181e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.389742803e+00 lpclm = -3.002097506e-07 wpclm = -6.253166196e-07 ppclm = 1.630738200e-13
+ pdiblc1 = 3.569721483e-01 lpdiblc1 = 3.176248153e-16 wpdiblc1 = 1.218537271e-15 ppdiblc1 = -2.324798132e-22
+ pdiblc2 = 8.406112145e-03 lpdiblc2 = -8.516243266e-18 wpdiblc2 = -3.267175419e-17 ppdiblc2 = 6.233315947e-24
+ pdiblcb = -1.032957699e-01 lpdiblcb = -2.521605147e-17 wpdiblcb = -9.673883916e-17 ppdiblcb = 1.845640307e-23
+ drout = 5.033266688e-01 ldrout = -1.682273876e-15 wdrout = -6.453880985e-15 pdrout = 1.231310165e-21
+ pscbe1 = 7.914198809e+08 lpscbe1 = -1.661944389e-07 wpscbe1 = -6.375885010e-07 ppscbe1 = 1.216430664e-13
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.662765292e-07 lalpha0 = -3.772961370e-14 walpha0 = -1.058933814e-13 palpha0 = 2.761551162e-20
+ alpha1 = 0.85
+ beta0 = 1.123895178e+01 lbeta0 = 8.034942409e-07 wbeta0 = 2.733891654e-06 pbeta0 = -7.129606690e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.003724933e-02 lkt1 = -4.196659342e-08 wkt1 = -1.177850524e-07 pkt1 = 3.071669265e-14
+ kt2 = -2.887893895e-02 lkt2 = -1.008054751e-17 wkt2 = -3.867306475e-17 pkt2 = 7.378278544e-24
+ at = -1.790597490e+05 lat = 5.418617662e-02 wat = 8.824448777e-02 pat = -2.301292699e-8
+ ute = -1.262490799e+00 lute = -1.474807435e-08 wute = -4.139251161e-08 pute = 1.079458756e-14
+ ua1 = -2.384732603e-11 lua1 = -1.902030267e-24 wua1 = -7.296954800e-24 pua1 = 1.392156823e-30
+ ub1 = 7.077531842e-19 lub1 = -2.701925638e-33 wub1 = -1.036567544e-32 pub1 = 1.977626141e-39
+ uc1 = 1.471862498e-10 luc1 = 3.912212746e-26 wuc1 = 1.500877862e-25 puc1 = -2.863471806e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.80 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {-7.924619035e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.178514156e-07 wvth0 = 9.400459055e-07 pvth0 = -1.516194797e-13
+ k1 = 0.90707349
+ k2 = -4.083638064e-01 lk2 = 4.388389027e-08 wk2 = 1.967510936e-07 pk2 = -3.344771707e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.584000555e-01 ldsub = 3.697184834e-11 wdsub = 1.453092562e-10 pdsub = -2.336369407e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999992e-03 lcdscd = 1.230168745e-18 wcdscd = 5.660125146e-18 pcdscd = -9.003995466e-25
+ cit = 0.0
+ voff = {-2.075299989e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.721580656e-16 wvoff = -7.836993277e-16 pvoff = 1.260079818e-22
+ nfactor = -6.537596072e+01 lnfactor = 1.091943640e-05 wnfactor = 4.223226157e-05 pnfactor = -6.843847262e-12
+ eta0 = 3.231038961e-02 leta0 = -5.195057784e-09 weta0 = -2.041796604e-08 peta0 = 3.282923088e-15
+ etab = -0.043998
+ u0 = -2.740290011e-02 lu0 = 9.830077904e-09 wu0 = 2.740134182e-08 pu0 = -5.012674006e-15
+ ua = 2.095541840e-09 lua = -5.605204870e-16 wua = -1.871097821e-15 pua = 3.268000561e-22
+ ub = -1.273520232e-17 lub = 2.635736298e-24 wub = 7.869843871e-24 pub = -1.460018959e-30
+ uc = 1.621727993e-09 luc = -2.483699919e-16 wuc = -9.761605222e-16 puc = 1.569529457e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.655766123e+06 lvsat = 4.744974360e-01 wvsat = 2.004571333e+00 pvsat = -3.271531937e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.132305965e-06 lb0 = -9.604577340e-13 wb0 = -2.854800955e-12 pb0 = 5.309583927e-19
+ b1 = -3.515314392e-06 lb1 = 6.578545512e-13 wb1 = 1.955363265e-12 pb1 = -3.636738702e-19
+ keta = -5.855695136e-01 lketa = 8.981015782e-08 wketa = 3.529779498e-07 pketa = -5.675391264e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.072893516e+00 lpclm = 1.696267822e-07 wpclm = 8.863854464e-07 ppclm = -1.253377703e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.609986601e-07 lalpha0 = 6.286711056e-14 walpha0 = 2.470845653e-13 palpha0 = -3.972773891e-20
+ alpha1 = 0.85
+ beta0 = 2.005574672e+01 lbeta0 = -8.786267981e-07 wbeta0 = -4.256155829e-06 pbeta0 = 6.206425301e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.739035193e-01 lkt1 = 3.317757676e-08 wkt1 = 1.704982743e-07 pkt1 = -2.428373011e-14
+ kt2 = -0.028878939
+ at = 3.795527042e+05 lat = -5.238925888e-02 wat = -2.059038048e-01 pat = 3.310644915e-8
+ ute = -2.444085418e+00 lute = 2.106836366e-07 wute = 6.273137034e-07 pute = -1.167851964e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.81 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.82 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.225219353e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.173473807e-06 wvth0 = 1.755577392e-08 pvth0 = -3.513048351e-13
+ k1 = 7.428610218e-01 lk1 = -3.498952003e-06 wk1 = -7.063348909e-08 pk1 = 1.413431635e-12
+ k2 = -1.089747373e-01 lk2 = 1.541600763e-06 wk2 = 3.443857457e-08 pk2 = -6.891429458e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.334255931e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.032263052e-07 wvoff = 1.721609947e-08 pvoff = -3.445076822e-13
+ nfactor = 4.723261510e+00 lnfactor = -1.602987046e-05 wnfactor = -1.981349644e-07 pnfactor = 3.964836372e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.021888796e-02 lu0 = 2.358353582e-07 wu0 = 5.042788863e-09 pu0 = -1.009101688e-13
+ ua = -1.738043863e-09 lua = 1.378540172e-14 wua = 2.713846733e-16 pua = -5.430620621e-21
+ ub = 1.361365732e-18 lub = -2.261533625e-24 wub = -3.731541830e-26 pub = 7.467108501e-31
+ uc = 6.580234079e-11 luc = -3.454930397e-16 wuc = -1.318359571e-18 puc = 2.638141124e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.160292432e+00 la0 = 4.048333449e-06 wa0 = 1.250485645e-07 pa0 = -2.502320063e-12
+ ags = 4.724837131e-01 lags = -2.553450595e-06 wags = -8.222347004e-08 pags = 1.645356263e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.630435158e-08 lb0 = 1.640891487e-12 wb0 = 4.578441793e-14 pb0 = -9.161821893e-19
+ b1 = 4.155395972e-08 lb1 = -5.838939187e-13 wb1 = -1.321865036e-14 pb1 = 2.645155835e-19
+ keta = -3.007770829e-02 lketa = 5.108975443e-07 wketa = 1.486276997e-08 pketa = -2.974157093e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.347719931e-01 lpclm = 3.034575526e-06 wpclm = 6.771135399e-08 ppclm = -1.354957415e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -6.833560397e-03 lpdiblc2 = 1.559618220e-07 wpdiblc2 = 4.001323413e-09 ppdiblc2 = -8.006962654e-14
+ pdiblcb = 1.025680820e+01 lpdiblcb = -2.057470637e-04 wpdiblcb = -5.572040884e-06 ppdiblcb = 1.115009177e-10
+ drout = 0.56
+ pscbe1 = -4.809228255e+08 lpscbe1 = 1.412607059e+04 wpscbe1 = 2.197636565e+02 ppscbe1 = -4.397643502e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.769214211e-01 lkt1 = -1.892735985e-07 wkt1 = -3.403857081e-09 pkt1 = 6.811385562e-14
+ kt2 = -3.518413649e-02 lkt2 = 1.133852255e-07 wkt2 = -1.659634346e-10 pkt2 = 3.321058774e-15
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -9.095327154e-01 lute = -4.119566177e-06 wute = -5.740833584e-08 pute = 1.148785923e-12
+ ua1 = 5.818406794e-10 lua1 = 1.078900178e-14 wua1 = 2.425883218e-16 pua1 = -4.854382994e-21
+ ub1 = 4.726390747e-20 lub1 = -1.234133024e-23 wub1 = -2.325545640e-25 pub1 = 4.653599614e-30
+ uc1 = 9.210253818e-11 luc1 = -1.166312177e-15 wuc1 = -1.226835950e-17 puc1 = 2.454995166e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.83 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.011796457e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.577148786e-07 wvth0 = -5.314882753e-08 pvth0 = 2.150945964e-13
+ k1 = 5.792489871e-01 lk1 = -2.188291007e-06 wk1 = -7.742138855e-08 pk1 = 1.467808045e-12
+ k2 = -4.773521515e-02 lk2 = 1.051024056e-06 wk2 = 3.720601738e-08 pk2 = -7.113123380e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.098697167e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.145252203e-07 wvoff = -4.404189257e-09 pvoff = -1.713121760e-13
+ nfactor = 3.087241344e-01 lnfactor = 1.933404375e-05 wnfactor = 1.997488264e-06 pnfactor = -1.362383145e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.463195597e-02 lu0 = -1.199482252e-07 wu0 = -1.675602394e-08 pu0 = 7.371545566e-14
+ ua = 1.499634463e-09 lua = -1.215094648e-14 wua = -1.340825671e-15 pua = 7.484451432e-21
+ ub = -1.239628140e-20 lub = 8.743379878e-24 wub = 7.394299124e-25 pub = -5.475629771e-30
+ uc = 1.271930437e-10 luc = -8.372808228e-16 wuc = -6.380674640e-17 puc = 5.269625056e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.049635017e+00 la0 = -3.075999680e-06 wa0 = -3.465071653e-07 pa0 = 1.275211975e-12
+ ags = 3.423043678e-01 lags = -1.510611718e-06 wags = 1.002101137e-08 pags = 9.064054629e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.785793739e-09 lb0 = 8.070476086e-13 wb0 = -4.920092209e-15 pb0 = -5.099992094e-19
+ b1 = -3.667485703e-08 lb1 = 4.278039133e-14 wb1 = 2.317601575e-14 pb1 = -2.703429826e-20
+ keta = 1.541054804e-02 lketa = 1.465008573e-07 wketa = -1.786332004e-08 pketa = -3.525400558e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.642642992e+00 lpclm = -1.120391555e-05 wpclm = -1.270153882e-06 ppclm = 9.362394691e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 3.081681516e-02 lpdiblc2 = -1.456472794e-07 wpdiblc2 = -1.760640615e-08 ppdiblc2 = 9.302527093e-14
+ pdiblcb = -3.087042461e+01 lpdiblcb = 1.237143972e-04 wpdiblcb = 1.671612265e-05 ppdiblcb = -6.704479071e-11
+ drout = 0.56
+ pscbe1 = 1.615700996e+09 lpscbe1 = -2.669534166e+03 wpscbe1 = -5.294692710e+02 ppscbe1 = 1.604301145e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.214738207e-01 lkt1 = 1.676261404e-07 wkt1 = 1.910149537e-08 pkt1 = -1.121717067e-13
+ kt2 = -8.604929512e-02 lkt2 = 5.208551261e-07 wkt2 = 4.137545168e-08 pkt2 = -3.294583278e-13
+ at = 140000.0
+ ute = -3.054447269e+00 lute = 1.306288530e-05 wute = 9.883429350e-07 pute = -7.228503717e-12
+ ua1 = -3.546451147e-10 lua1 = 1.829098907e-14 wua1 = 1.014927243e-15 pua1 = -1.104142481e-20
+ ub1 = -3.748327798e-19 lub1 = -8.960004008e-24 wub1 = -3.545141521e-25 pub1 = 5.630591775e-30
+ uc1 = 2.169604830e-10 luc1 = -2.166522453e-15 wuc1 = -1.564087500e-16 puc1 = 1.400177339e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.84 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {3.170859599e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.817240990e-07 wvth0 = 1.222905854e-07 pvth0 = -4.885553449e-13
+ k1 = -2.709787118e-01 lk1 = 1.221790345e-06 wk1 = 4.498077842e-07 pk1 = -6.467953404e-13
+ k2 = 4.031671796e-01 lk2 = -7.574489557e-07 wk2 = -2.430005125e-07 pk2 = 4.125360891e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.256182131e+00 ldsub = 7.284317864e-06 wdsub = 1.147703606e-06 pdsub = -4.603193557e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {2.240673878e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.024825043e-06 wvoff = -1.959827088e-07 pvoff = 5.970682679e-13
+ nfactor = 1.364038402e+01 lnfactor = -3.413639107e-05 wnfactor = -6.376575489e-06 pnfactor = 1.996274622e-11
+ eta0 = -4.012882647e-01 leta0 = 1.930344234e-06 weta0 = 3.041414557e-07 peta0 = -1.219846292e-12
+ etab = 3.507488603e-01 letab = -1.687533639e-06 wetab = -2.658846688e-07 petab = 1.066406507e-12
+ u0 = 2.806354577e-02 lu0 = -1.338801750e-08 wu0 = 8.038198033e-10 pu0 = 3.286680199e-15
+ ua = 2.557894949e-09 lua = -1.639540283e-14 wua = -1.769021654e-15 pua = 9.201853888e-21
+ ub = -4.302580468e-18 lub = 2.595039055e-23 wub = 3.135343290e-24 pub = -1.508512560e-29
+ uc = -2.379563201e-10 luc = 6.272551334e-16 wuc = 1.481636926e-16 puc = -3.232055636e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 9.028145105e-01 la0 = 1.523651952e-06 wa0 = 3.871902937e-07 pa0 = -1.667491522e-12
+ ags = -1.000395022e+00 lags = 3.874668198e-06 wags = 7.185362784e-07 pags = -1.935297651e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.042275371e-07 lb0 = -3.819167856e-13 wb0 = -1.922511160e-13 pb0 = 2.413454382e-19
+ b1 = 4.089175861e-08 lb1 = -2.683227047e-13 wb1 = -2.584081080e-14 pb1 = 1.695617035e-19
+ keta = 1.969736027e-01 lketa = -5.817097006e-07 wketa = -1.064868830e-07 pketa = 3.201961399e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.179382640e+00 lpclm = 8.136197346e-06 wpclm = 2.330870809e-06 ppclm = -5.080544728e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -4.948768676e-03 lpdiblc2 = -2.199176451e-09 wpdiblc2 = 4.000513243e-09 ppdiblc2 = 6.364541126e-15
+ pdiblcb = 5.067425545e-02 lpdiblcb = -3.035132443e-07 wpdiblcb = -4.782098360e-08 ppdiblcb = 1.917997315e-13
+ drout = 0.56
+ pscbe1 = 1.101033985e+09 lpscbe1 = -6.053149235e+02 wpscbe1 = -2.596433974e+02 ppscbe1 = 5.220873084e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.227282992e-01 lkt1 = 9.748147854e-07 wkt1 = 1.434342517e-07 pkt1 = -6.108437850e-13
+ kt2 = -7.938462818e-02 lkt2 = 4.941245733e-07 wkt2 = 3.517995610e-08 pkt2 = -3.046095209e-13
+ at = 1.578766074e+05 lat = -7.169924669e-02 wat = 7.000991999e-03 pat = -2.807948069e-8
+ ute = -7.087306456e+00 lute = 2.923782047e-05 wute = 3.371484071e-06 pute = -1.678677282e-11
+ ua1 = -1.800301168e-08 lua1 = 8.907481063e-14 wua1 = 1.092717142e-14 pua1 = -5.079731497e-20
+ ub1 = 1.499778034e-17 lub1 = -7.061626550e-23 wub1 = -8.940876022e-24 pub1 = 4.006865175e-29
+ uc1 = -9.229235894e-11 luc1 = -9.261754840e-16 wuc1 = 5.435028445e-17 puc1 = 5.548679539e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.85 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {7.937800972e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.680579848e-08 wvth0 = -1.640195908e-07 pvth0 = 8.715314912e-14
+ k1 = 6.484758779e-01 lk1 = -6.270360717e-07 wk1 = -3.049074960e-08 pk1 = 3.189822272e-13
+ k2 = -1.005150039e-01 lk2 = 2.553481272e-07 wk2 = 3.104208571e-08 pk2 = -1.385049307e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.495600062e+00 ldsub = -4.281285244e-06 wdsub = -2.295407213e-06 pdsub = 2.320165475e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-3.198180790e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.881223899e-08 wvoff = 1.388585976e-07 pvoff = -7.622594312e-14
+ nfactor = -6.058513806e+00 lnfactor = 5.473876890e-06 wnfactor = 5.572404867e-06 pnfactor = -4.064096199e-12
+ eta0 = 1.120880502e+00 leta0 = -1.130411413e-06 weta0 = -6.082827191e-07 peta0 = 6.148434642e-13
+ etab = -8.969676719e-01 letab = 8.213572965e-07 wetab = 5.317693376e-07 petab = -5.375050017e-13
+ u0 = 1.602787924e-02 lu0 = 1.081313225e-08 wu0 = 7.487636141e-09 pu0 = -1.015304412e-14
+ ua = -8.248751638e-09 lua = 5.334450837e-15 wua = 4.632663562e-15 pua = -3.670565122e-21
+ ub = 1.230099358e-17 lub = -7.435843687e-24 wub = -6.825140103e-24 pub = 4.943274956e-30
+ uc = -1.083141739e-10 luc = 3.665725207e-16 wuc = 9.237901644e-17 puc = -2.110345177e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.981918887e+04 lvsat = 1.009028725e-01 wvsat = 2.532338016e-02 pvsat = -5.091989829e-8
+ a0 = 7.116585410e+00 la0 = -1.097091158e-05 wa0 = -3.593451700e-06 pa0 = 6.336727671e-12
+ ags = 4.409992822e+00 lags = -7.004463935e-06 wags = -2.555445842e-06 pags = 4.647979762e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.401602900e-07 lb0 = -4.541698620e-13 wb0 = -2.149581724e-13 pb0 = 2.870044692e-19
+ b1 = 7.060957997e-10 lb1 = -1.875179366e-13 wb1 = -4.462045309e-16 pb1 = 1.184985847e-19
+ keta = -6.348267072e-01 lketa = 1.090862717e-06 wketa = 3.838371632e-07 pketa = -6.657405877e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.155315110e+00 lpclm = -2.590738205e-06 wpclm = -1.093786105e-06 ppclm = 1.805707450e-12
+ pdiblc1 = 5.371846616e-01 lpdiblc1 = -2.959568570e-07 wpdiblc1 = -6.024587525e-08 ppdiblc1 = 1.211415625e-13
+ pdiblc2 = -2.478774381e-02 lpdiblc2 = 3.769275700e-08 wpdiblc2 = 1.868584952e-08 ppdiblc2 = -2.316452746e-14
+ pdiblcb = 1.476230808e-01 lpdiblcb = -4.984565851e-07 wpdiblcb = -9.351813708e-08 ppdiblcb = 2.836869280e-13
+ drout = 3.904020436e+00 ldrout = -6.724109477e-06 wdrout = -2.009269098e-06 pdrout = 4.040210173e-12
+ pscbe1 = 3.976706747e+08 lpscbe1 = 8.089981747e+02 wpscbe1 = 2.542447752e+02 ppscbe1 = -5.112318345e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.345293063e-05 lalpha0 = -6.720636099e-11 walpha0 = -2.112025290e-11 palpha0 = 4.246830885e-17
+ alpha1 = 1.935871632e+00 lalpha1 = -2.183455474e-06 walpha1 = -5.884685850e-07 palpha1 = 1.183284392e-12
+ beta0 = 3.579543680e+01 lbeta0 = -4.410746922e-05 wbeta0 = -1.386170445e-05 pbeta0 = 2.787292124e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 7.346911206e-02 lkt1 = -2.240106225e-07 wkt1 = -2.531311393e-07 pkt1 = 1.865643512e-13
+ kt2 = 4.265088998e-01 lkt2 = -5.231190502e-07 wkt2 = -2.688742999e-07 pkt2 = 3.067785203e-13
+ at = 1.896562588e+04 lat = 2.076210102e-01 wat = 7.456434576e-02 pat = -1.639349266e-7
+ ute = 1.587559330e+01 lute = -1.693565688e-05 wute = -9.900478187e-06 pute = 9.900303079e-12
+ ua1 = 5.182949306e-08 lua1 = -5.134341226e-14 wua1 = -2.896074252e-14 pua1 = 2.940874395e-20
+ ub1 = -3.909037288e-17 lub1 = 3.814343576e-23 wub1 = 2.171600247e-23 pub1 = -2.157577033e-29
+ uc1 = -9.901999276e-10 luc1 = 8.793244844e-16 wuc1 = 5.758124179e-16 puc1 = -4.936808036e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.86 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {8.424746912e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.260256124e-07 wvth0 = -1.572711140e-07 pvth0 = 8.033188323e-14
+ k1 = -4.283618718e-01 lk1 = 4.614164500e-07 wk1 = 5.763252088e-07 pk1 = -2.943788481e-13
+ k2 = 3.152370518e-01 lk2 = -1.648882301e-07 wk2 = -2.142560502e-07 pk2 = 1.094389909e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667334e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-3.621758405e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.116268713e-07 wvoff = 1.282607666e-07 pvoff = -6.551380394e-14
+ nfactor = -4.171259751e+00 lnfactor = 3.566266913e-06 wnfactor = 3.136825254e-06 pnfactor = -1.602246424e-12
+ eta0 = -4.954524662e-01 leta0 = 5.033553234e-07 weta0 = -3.846199902e-13 peta0 = 1.964585063e-19
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 3.501386970e-02 lu0 = -8.377641105e-09 wu0 = -5.169292668e-09 pu0 = 2.640402325e-15
+ ua = -4.378955446e-09 lua = 1.422915023e-15 wua = 2.024132699e-15 pua = -1.033898645e-21
+ ub = 8.328205928e-18 lub = -3.420205550e-24 wub = -3.910962216e-24 pub = 1.997664746e-30
+ uc = 4.605098122e-10 luc = -2.083868008e-16 wuc = -2.353182024e-16 puc = 1.201972433e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.317214727e+05 lvsat = 2.641859117e-01 wvsat = -5.064676031e-02 pvsat = 2.586965611e-8
+ a0 = -8.969601952e+00 la0 = 5.288781398e-06 wa0 = 5.409034001e-06 pa0 = -2.762858841e-12
+ ags = -5.253430486e+00 lags = 2.763189057e-06 wags = 4.129941761e-06 pags = -2.109516432e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.206812063e-07 lb0 = 1.127208706e-13 wb0 = 1.394555161e-13 pb0 = -7.123192522e-20
+ b1 = -3.736084496e-07 lb1 = 1.908339655e-13 wb1 = 2.360951348e-13 pb1 = -1.205940895e-19
+ keta = 9.056443002e-01 lketa = -4.662238103e-07 wketa = -5.555267136e-07 pketa = 2.837552680e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.285908178e+00 lpclm = 8.876021169e-07 wpclm = 1.400247536e-06 ppclm = -7.152268381e-13
+ pdiblc1 = 4.602994019e-01 lpdiblc1 = -2.182423128e-07 wpdiblc1 = 1.204917505e-07 ppdiblc1 = -6.154549928e-14
+ pdiblc2 = 2.522786576e-02 lpdiblc2 = -1.286232093e-08 wpdiblc2 = -8.554264740e-09 ppdiblc2 = 4.369398669e-15
+ pdiblcb = -6.018364499e-01 lpdiblcb = 2.590866161e-07 wpdiblcb = 3.783202085e-07 ppdiblcb = -1.932406660e-13
+ drout = -6.577532450e+00 ldrout = 3.870497439e-06 wdrout = 4.018538197e-06 pdrout = -2.052613051e-12
+ pscbe1 = 1.975543419e+09 lpscbe1 = -7.858935053e+02 wpscbe1 = -5.084895504e+02 ppscbe1 = 2.597293435e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -7.076934490e-05 lalpha0 = 3.814005601e-11 walpha0 = 4.224050580e-11 palpha0 = -2.157585900e-17
+ alpha1 = -1.321743263e+00 lalpha1 = 1.109296054e-06 walpha1 = 1.176937170e-06 palpha1 = -6.011630293e-13
+ beta0 = -3.425856997e+01 lbeta0 = 2.670214007e-05 wbeta0 = 2.772340889e-05 pbeta0 = -1.416072914e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.453106478e-02 lkt1 = -1.350612757e-07 wkt1 = -1.385941211e-07 pkt1 = 7.079193675e-14
+ kt2 = -1.465089572e-01 lkt2 = 5.607937740e-08 wkt2 = 7.000828446e-08 pkt2 = -3.575925159e-14
+ at = 4.426972833e+05 lat = -2.206810169e-01 wat = -1.771326595e-01 pat = 9.047688263e-8
+ ute = -4.391146268e-01 lute = -4.449785145e-07 wute = -2.139233308e-07 pute = 1.092690425e-13
+ ua1 = 1.240617085e-09 lua1 = -2.088846656e-16 wua1 = 2.712617097e-16 pua1 = -1.385566837e-22
+ ub1 = -2.091621868e-18 lub1 = 7.456162207e-25 wub1 = 7.489218910e-25 pub1 = -3.825388170e-31
+ uc1 = -2.489757399e-10 luc1 = 1.301054526e-16 wuc1 = 1.766846542e-16 puc1 = -9.024804776e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.87 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.375477052e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.135177687e-8
+ k1 = 2.425254328e-02 lk1 = 2.302273434e-7
+ k2 = 1.380233204e-01 lk2 = -7.436993714e-08 wk2 = 6.938893904e-24 pk2 = 8.673617380e-30
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988867e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
+ voff = {-1.072895691e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.856546770e-8
+ nfactor = 4.181852128e+00 lnfactor = -7.003856916e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928473e-02 letab = -2.311014722e-08 wetab = 7.806255642e-24 petab = 6.288372600e-30
+ u0 = 1.686628126e-02 lu0 = 8.918930054e-10
+ ua = -2.102030833e-09 lua = 2.598938077e-16
+ ub = 2.286030910e-18 lub = -3.339471417e-25 wub = -1.540743956e-39
+ uc = 1.078724766e-11 luc = 2.132518900e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.032128435e+05 lvsat = -6.012964798e-2
+ a0 = 1.264221183e+00 la0 = 6.148781439e-8
+ ags = -9.846887479e-01 lags = 5.827755398e-07 wags = 2.220446049e-22 pags = -1.110223025e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.684190351e-18 lb0 = 1.221571265e-24
+ b1 = -2.709394687e-17 lb1 = 7.065722030e-24
+ keta = 7.220181439e-02 lketa = -4.051305669e-08 wketa = 1.387778781e-23 pketa = -3.469446952e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500260e-01 lpclm = -1.136192512e-07 wpclm = 4.440892099e-22
+ pdiblc1 = -3.048846467e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = -1.110223025e-22 ppdiblc1 = 1.387778781e-29
+ pdiblc2 = -8.673906562e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 1.084202172e-25 ppdiblc2 = 5.692061406e-31
+ pdiblcb = -8.553970445e-02 lpdiblcb = -4.630533311e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076329e+07 lpscbe1 = 1.888714223e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729690e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380752e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373076e+03 lat = 9.625574770e-03 pat = 3.637978807e-24
+ ute = -1.301136473e+00 lute = -4.669823644e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393852e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873018e-25 wub1 = -7.703719778e-40
+ uc1 = -1.418079324e-10 luc1 = 7.536563684e-17 wuc1 = 4.523643975e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.88 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.910376278e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610889862e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456657017e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
+ voff = {-9.930380979e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149736110e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935927057e-16
+ ags = 1.250000000e+00 lags = 6.286171583e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026246086e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347658096e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990252573e-18
+ drout = 5.033266586e-01 ldrout = 2.662110532e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629947662e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595196197e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009865455e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275664625e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190826499e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.89 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {1.140963279e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.071407151e-07 wvth0 = -2.817473370e-07 pvth0 = 5.375344743e-14
+ k1 = 0.90707349
+ k2 = -1.379104027e-02 lk2 = -2.492342843e-08 wk2 = -5.259206361e-08 pk2 = 1.003382945e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999998e-03 lcdscd = 4.335403564e-19 wcdscd = 2.080779993e-18 pcdscd = -3.969845286e-25
+ cit = 0.0
+ voff = {-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.724287462e-17
+ nfactor = -1.367122711e+00 lnfactor = 6.277113832e-07 wnfactor = 1.783028553e-06 pnfactor = -3.401768854e-13
+ eta0 = 1.642889168e-09 leta0 = -2.641230358e-16 weta0 = 5.415415969e-19 peta0 = -1.033185551e-25
+ etab = -0.043998
+ u0 = -1.317993572e-01 lu0 = 3.008787420e-08 wu0 = 9.337280374e-08 pu0 = -1.781422373e-14
+ ua = 5.036359176e-10 lua = -3.045641810e-16 wua = -8.651215275e-16 pua = 1.650530758e-22
+ ub = -1.054947243e-17 lub = 2.284301680e-24 wub = 6.488611209e-24 pub = -1.237936178e-30
+ uc = 7.700399983e-11 luc = 2.675329576e-26 wuc = -1.431022460e-28 puc = 2.724526143e-35
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.500760136e+06 lvsat = -4.218004844e-01 wvsat = -1.254002619e+00 pvsat = 2.392461438e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.409772263e-06 lb0 = -8.442842676e-13 wb0 = -2.398208787e-12 pb0 = 4.575446617e-19
+ b1 = -3.020423958e-06 lb1 = 5.782830229e-13 wb1 = 1.642626163e-12 pb1 = -3.133900752e-19
+ keta = -2.700000009e-02 lketa = 1.436820107e-17 wketa = 8.160139231e-20 pketa = -1.557087792e-26
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.236013226e+00 lpclm = -2.016130945e-07 wpclm = -5.726866092e-07 ppclm = 1.092605874e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.200778689e-24 walpha0 = -1.631597215e-25 palpha0 = 3.112846081e-32
+ alpha1 = 0.85
+ beta0 = 1.005373824e+01 lbeta0 = 7.267793524e-07 wbeta0 = 2.064433393e-06 pbeta0 = -3.938649894e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.839584507e-02 lkt1 = -3.686397382e-08 wkt1 = -1.047129613e-07 pkt1 = 1.997776703e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.577747753e-11 wat = -3.469176590e-14 pat = 6.635673344e-21
+ ute = -2.268108645e+00 lute = 1.816948390e-07 wute = 5.161083492e-07 pute = -9.846624750e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.90 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.91 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.549167264e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016575863e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-07 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = -1.525878906e-17
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-08 wkt1 = -1.776356839e-21
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16 puc1 = -1.654361225e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.92 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.031067740e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179965467e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647566e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-08 wketa = -5.551115123e-23 pketa = -2.220446049e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = -4.440892099e-22 ppclm = -3.552713679e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267872e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.93 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.427426575e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.375696972e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15 wua1 = -6.617444900e-30 pua1 = -1.323488980e-35
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.94 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.911229542e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.358925766e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159063e-03 leta0 = 4.128463499e-09 weta0 = 3.469446952e-24 peta0 = 3.469446952e-30
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -1.561251128e-22 petab = -2.949029909e-28
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = 1.665334537e-22 pketa = -5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 5.929230631e-27 palpha0 = 1.312901068e-32
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -1.654361225e-30 pua1 = 4.963083675e-36
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 pub1 = -1.540743956e-45
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17 wuc1 = 4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.95 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.522701748e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.220679177e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610700e-8
+ k2 = -8.011891576e-02 lk2 = 3.705406310e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667334e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.255026663e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.262472634e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217668e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -2.498001805e-22 peta0 = -6.938893904e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.547523263e-02 lu0 = -3.505438827e-9
+ ua = -6.439246683e-10 lua = -4.848864078e-16
+ ub = 1.111503064e-18 lub = 2.659852385e-25
+ uc = 2.628890916e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.251774050e+05 lvsat = 3.119218935e-1
+ a0 = 1.011417809e+00 la0 = 1.906162389e-7
+ ags = 2.367344374e+00 lags = -1.129396050e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608784e-08 lb1 = -3.169227303e-14
+ keta = -1.194413445e-01 lketa = 5.737558588e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701757e-07 wpclm = 7.105427358e-21
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109111e-03 lpdiblc2 = -4.799688221e-9
+ pdiblcb = 9.625889888e-02 lpdiblcb = -9.749071472e-08 wpdiblcb = -1.422473250e-22 ppdiblcb = 1.066854938e-28
+ drout = 8.376749865e-01 ldrout = 8.291329324e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279453e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552323e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457427e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380072e-9
+ at = 1.158432509e+05 lat = -5.372855309e-2
+ ute = -8.338566439e-01 lute = -2.433498185e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563802e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648484e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475370e-17 wuc1 = 4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.96 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.375477052e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.135177687e-8
+ k1 = 2.425254328e-02 lk1 = 2.302273434e-7
+ k2 = 1.380233204e-01 lk2 = -7.436993714e-08 wk2 = -2.220446049e-22 pk2 = 5.551115123e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988867e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-09 wcdscd = 5.551115123e-23
+ cit = 0.0
+ voff = {-1.072895691e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.856546770e-8
+ nfactor = 4.181852128e+00 lnfactor = -7.003856916e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928473e-02 letab = -2.311014722e-08 wetab = 1.387778781e-23 petab = -5.204170428e-29
+ u0 = 1.686628126e-02 lu0 = 8.918930054e-10
+ ua = -2.102030833e-09 lua = 2.598938077e-16 wua = 1.323488980e-29
+ ub = 2.286030910e-18 lub = -3.339471417e-25
+ uc = 1.078724766e-11 luc = 2.132518900e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.032128435e+05 lvsat = -6.012964798e-2
+ a0 = 1.264221183e+00 la0 = 6.148781439e-8
+ ags = -9.846887479e-01 lags = 5.827755398e-07 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.684190351e-18 lb0 = 1.221571265e-24
+ b1 = -2.709394687e-17 lb1 = 7.065722030e-24
+ keta = 7.220181439e-02 lketa = -4.051305669e-08 wketa = -5.551115123e-23 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500260e-01 lpclm = -1.136192512e-7
+ pdiblc1 = -3.048846467e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = 2.220446049e-22 ppdiblc1 = -4.440892099e-28
+ pdiblc2 = -8.673906562e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 2.125036258e-23 ppdiblc2 = 2.385244779e-30
+ pdiblcb = -8.553970445e-02 lpdiblcb = -4.630533311e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076329e+07 lpscbe1 = 1.888714223e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729690e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380752e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373076e+03 lat = 9.625574770e-03 pat = 2.910383046e-23
+ ute = -1.301136473e+00 lute = -4.669823644e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393852e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873018e-25 pub1 = 1.540743956e-45
+ uc1 = -1.418079324e-10 luc1 = 7.536563684e-17 wuc1 = -5.169878828e-32 puc1 = 1.421716678e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.97 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.910376278e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456612608e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
+ voff = {-9.930380979e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149569577e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.936033638e-16
+ ags = 1.250000000e+00 lags = 6.285461041e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026379313e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347644218e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990141551e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629852295e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009866231e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190619704e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.98 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {-3.567178047e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.911067358e-07 wvth0 = 2.269745108e-06 pvth0 = -4.330355901e-13
+ k1 = 0.90707349
+ k2 = -1.802308111e+00 lk2 = 3.163005895e-07 wk2 = 9.166625698e-07 pk2 = -1.748863850e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000027e-03 lcdscd = -5.141442827e-18 wcdscd = -1.375510816e-17 pcdscd = 2.624282736e-24
+ cit = 0.0
+ voff = {-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.724220849e-17
+ nfactor = -1.367121211e+00 lnfactor = 6.277110970e-07 wnfactor = 1.783027739e-06 pnfactor = -3.401767303e-13
+ eta0 = 1.642889326e-09 leta0 = -2.641230346e-16 weta0 = 5.415449217e-19 peta0 = -1.033191894e-25
+ etab = -0.043998
+ u0 = 1.025634817e+00 lu0 = -1.907343621e-07 wu0 = -5.338778131e-07 pu0 = 1.018564124e-13
+ ua = 5.036486647e-10 lua = -3.045666130e-16 wua = -8.651284356e-16 pua = 1.650543937e-22
+ ub = -1.054935338e-17 lub = 2.284278967e-24 wub = 6.488546693e-24 pub = -1.237923869e-30
+ uc = 7.700399983e-11 luc = 2.713483281e-26 wuc = 9.429858983e-28 puc = -1.799117832e-34
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.989946961e+07 lvsat = 3.851849748e+00 wvsat = 1.088539869e+01 pvsat = -2.076781674e-6
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.409769924e-06 lb0 = -8.442838214e-13 wb0 = -2.398207520e-12 pb0 = 4.575444199e-19
+ b1 = -3.020424216e-06 lb1 = 5.782830722e-13 wb1 = 1.642626303e-12 pb1 = -3.133901019e-19
+ keta = -2.700000009e-02 lketa = 1.414912632e-17 wketa = -5.409006576e-19 pketa = 1.032507413e-25
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.236013822e+00 lpclm = -2.016132082e-07 wpclm = -5.726869319e-07 ppclm = 1.092606490e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -2.762597957e-24 walpha0 = 1.081661074e-24 palpha0 = -2.063584018e-31
+ alpha1 = 0.85
+ beta0 = 1.011879351e+01 lbeta0 = 7.143677172e-07 wbeta0 = 2.029177860e-06 pbeta0 = -3.871387271e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.440041678e-02 lkt1 = -3.571838560e-08 wkt1 = -1.014588917e-07 pkt1 = 1.935693611e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.587113366e-11 wat = 2.309679985e-13 pat = -4.423782229e-20
+ ute = -2.251844814e+00 lute = 1.785919276e-07 wute = 5.072944585e-07 pute = -9.678468056e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.99 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.100 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.549167264e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016575863e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14 wb1 = 2.646977960e-29
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-07 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = -3.814697266e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.101 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.031067740e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179965467e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647567e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = 4.440892099e-22 ppclm = 2.664535259e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-08 ppdiblc2 = -1.387778781e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267872e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.102 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.427426575e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.375696972e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-06 wpclm = 1.776356839e-21
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.103 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.911229542e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.358925766e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159062e-03 leta0 = 4.128463499e-09 peta0 = -3.469446952e-30
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = 1.734723476e-24 petab = -4.510281038e-29
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24
+ uc = 6.214820228e-11 luc = -2.283891413e-17 wuc = 1.033975766e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 pb0 = -5.293955920e-35
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = 1.387778781e-23 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = -7.411538288e-28 palpha0 = -1.799945013e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-02 wat = 2.328306437e-16
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -8.271806126e-31
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 pub1 = 7.703719778e-46
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.104 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.522701748e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.220679177e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610700e-8
+ k2 = -8.011891576e-02 lk2 = 3.705406310e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667334e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.255026663e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.262472634e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217668e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -4.024558464e-22 peta0 = -2.775557562e-29
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.547523263e-02 lu0 = -3.505438827e-9
+ ua = -6.439246683e-10 lua = -4.848864078e-16
+ ub = 1.111503064e-18 lub = 2.659852385e-25
+ uc = 2.628890916e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.251774050e+05 lvsat = 3.119218935e-1
+ a0 = 1.011417809e+00 la0 = 1.906162389e-7
+ ags = 2.367344374e+00 lags = -1.129396050e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608784e-08 lb1 = -3.169227303e-14
+ keta = -1.194413445e-01 lketa = 5.737558588e-08 pketa = -1.110223025e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701757e-7
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109111e-03 lpdiblc2 = -4.799688221e-9
+ pdiblcb = 9.625889888e-02 lpdiblcb = -9.749071472e-08 wpdiblcb = -4.640385298e-23 ppdiblcb = 5.247538515e-29
+ drout = 8.376749865e-01 ldrout = 8.291329324e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279453e+02 wpscbe1 = 1.907348633e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552323e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457427e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380072e-9
+ at = 1.158432509e+05 lat = -5.372855309e-2
+ ute = -8.338566439e-01 lute = -2.433498185e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563802e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648484e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475370e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.105 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.375477052e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.135177687e-8
+ k1 = 2.425254328e-02 lk1 = 2.302273434e-7
+ k2 = 1.380233204e-01 lk2 = -7.436993714e-08 wk2 = -8.326672685e-23 pk2 = 3.469446952e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988867e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
+ voff = {-1.072895691e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.856546770e-8
+ nfactor = 4.181852128e+00 lnfactor = -7.003856916e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928473e-02 letab = -2.311014722e-08 wetab = 1.561251128e-23 petab = 9.540979118e-30
+ u0 = 1.686628126e-02 lu0 = 8.918930054e-10
+ ua = -2.102030833e-09 lua = 2.598938077e-16
+ ub = 2.286030910e-18 lub = -3.339471417e-25
+ uc = 1.078724766e-11 luc = 2.132518900e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.032128435e+05 lvsat = -6.012964798e-2
+ a0 = 1.264221183e+00 la0 = 6.148781439e-8
+ ags = -9.846887479e-01 lags = 5.827755398e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.684190351e-18 lb0 = 1.221571265e-24
+ b1 = -2.709394687e-17 lb1 = 7.065722030e-24
+ keta = 7.220181439e-02 lketa = -4.051305669e-08 wketa = -2.775557562e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500260e-01 lpclm = -1.136192512e-7
+ pdiblc1 = -3.048846467e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = -2.220446049e-22 ppdiblc1 = -8.326672685e-29
+ pdiblc2 = -8.673906562e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = -1.951563910e-24 ppdiblc2 = 1.219727444e-30
+ pdiblcb = -8.553970445e-02 lpdiblcb = -4.630533311e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076329e+07 lpscbe1 = 1.888714223e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729690e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380752e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373076e+03 lat = 9.625574770e-03 pat = 7.275957614e-24
+ ute = -1.301136473e+00 lute = -4.669823644e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393852e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873018e-25 wub1 = -1.540743956e-39 pub1 = -3.851859889e-46
+ uc1 = -1.418079324e-10 luc1 = 7.536563684e-17 wuc1 = -3.877409121e-32 puc1 = -6.462348536e-39
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.106 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.910376278e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610978680e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456701426e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
+ voff = {-9.930380979e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149680599e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935962584e-16
+ ags = 1.250000000e+00 lags = 6.286171583e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026290495e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347671974e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990141551e-18
+ drout = 5.033266586e-01 ldrout = 2.662110532e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629852295e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009864680e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190826499e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.107 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {1.625879187e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.996558816e-07 wvth0 = -4.926082127e-07 pvth0 = 9.398275046e-14
+ k1 = 0.90707349
+ k2 = 2.979877433e-01 lk2 = -8.440645544e-08 wk2 = -2.005520048e-07 pk2 = 3.826251479e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.584979911e-01 ldsub = 2.518544814e-11 wdsub = 7.021975303e-11 pdsub = -1.339694580e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079655892e-19
+ cit = 0.0
+ voff = {-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.724309667e-17
+ nfactor = 1.334758346e+01 lnfactor = -2.179648549e-06 wnfactor = -6.044194547e-06 pnfactor = 1.153147701e-12
+ eta0 = 1.826783307e-02 leta0 = -3.485246401e-09 weta0 = -9.717243132e-09 peta0 = 1.853913948e-15
+ etab = -0.043998
+ u0 = -3.317912352e-01 lu0 = 6.824352463e-08 wu0 = 1.881805416e-07 pu0 = -3.590221282e-14
+ ua = -3.087980150e-09 lua = 3.806658820e-16 wua = 1.045373863e-15 pua = -1.994426978e-22
+ ub = 2.653989546e-17 lub = -4.791830462e-24 wub = -1.324041162e-23 pub = 2.526085172e-30
+ uc = 3.575979994e-10 luc = -5.353340678e-17 wuc = -1.492569274e-16 puc = 2.847613215e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.124878107e+07 lvsat = -2.090800406e+00 wvsat = -5.683352593e+00 pvsat = 1.084304108e-6
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.325206324e-05 lb0 = 2.525346681e-12 wb0 = 6.996686721e-12 pb0 = -1.334869873e-18
+ b1 = 2.663302983e-06 lb1 = -5.060925053e-13 wb1 = -1.380730074e-12 pb1 = 2.634239678e-19
+ keta = -2.700000009e-02 lketa = 1.434302677e-17
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.564203824e-01 lpclm = 1.022009439e-07 wpclm = 2.743797791e-07 ppclm = -5.234782053e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.150539047e-24
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968377e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.983091395e-01 lkt1 = 5.088104398e-08 wkt1 = 1.399896830e-07 pkt1 = -2.670807166e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.578824595e-11
+ ute = 4.121252916e-01 lute = -3.296562729e-07 wute = -9.097564876e-07 pute = 1.735688012e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.108 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.109 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.549167264e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016575863e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.110 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.031067740e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179965467e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647566e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = 1.332267630e-21
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267871e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16 puc1 = -8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.111 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.427426575e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.375696972e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-01 wat = -9.313225746e-16
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.112 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.911229542e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.358925766e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159062e-03 leta0 = 4.128463499e-09 peta0 = -6.938893904e-30
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -1.873501354e-22 petab = 1.734723476e-28
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15 pua = -3.308722450e-36
+ ub = -2.930959084e-19 lub = 1.685734216e-24 pub = -3.081487911e-45
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = -2.775557562e-23 pketa = 2.220446049e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 7.623296525e-27 palpha0 = -6.988021815e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -1.654361225e-30
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 pub1 = 1.540743956e-45
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.113 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.522701748e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.220679177e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610700e-8
+ k2 = -8.011891576e-02 lk2 = 3.705406310e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667334e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.255026663e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.262472634e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217668e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 4.718447855e-22 peta0 = 6.245004514e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.547523263e-02 lu0 = -3.505438827e-9
+ ua = -6.439246683e-10 lua = -4.848864078e-16
+ ub = 1.111503064e-18 lub = 2.659852385e-25
+ uc = 2.628890916e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.251774050e+05 lvsat = 3.119218935e-01 wvsat = 4.656612873e-16 pvsat = -4.656612873e-22
+ a0 = 1.011417809e+00 la0 = 1.906162389e-7
+ ags = 2.367344374e+00 lags = -1.129396050e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608784e-08 lb1 = -3.169227303e-14
+ keta = -1.194413445e-01 lketa = 5.737558588e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701757e-07 wpclm = -7.105427358e-21
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109111e-03 lpdiblc2 = -4.799688221e-9
+ pdiblcb = 9.625889888e-02 lpdiblcb = -9.749071472e-08 wpdiblcb = -3.122502257e-23 ppdiblcb = 1.847480502e-28
+ drout = 8.376749865e-01 ldrout = 8.291329324e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279453e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552323e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457427e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380072e-9
+ at = 1.158432509e+05 lat = -5.372855309e-2
+ ute = -8.338566439e-01 lute = -2.433498185e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563802e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648484e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475370e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.114 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.375477052e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.135177687e-8
+ k1 = 2.425254328e-02 lk1 = 2.302273434e-7
+ k2 = 1.380233204e-01 lk2 = -7.436993714e-08 wk2 = 5.551115123e-23 pk2 = -8.326672685e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988867e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
+ voff = {-1.072895691e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.856546770e-8
+ nfactor = 4.181852128e+00 lnfactor = -7.003856916e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928473e-02 letab = -2.311014722e-08 wetab = 2.775557562e-23 petab = -3.816391647e-29
+ u0 = 1.686628126e-02 lu0 = 8.918930054e-10
+ ua = -2.102030833e-09 lua = 2.598938077e-16
+ ub = 2.286030910e-18 lub = -3.339471417e-25
+ uc = 1.078724766e-11 luc = 2.132518900e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.032128435e+05 lvsat = -6.012964798e-2
+ a0 = 1.264221183e+00 la0 = 6.148781439e-8
+ ags = -9.846887479e-01 lags = 5.827755398e-07 wags = 1.776356839e-21 pags = 8.881784197e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.684190351e-18 lb0 = 1.221571265e-24
+ b1 = -2.709394687e-17 lb1 = 7.065722030e-24
+ keta = 7.220181439e-02 lketa = -4.051305669e-08 wketa = -1.110223025e-22 pketa = -1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500260e-01 lpclm = -1.136192512e-7
+ pdiblc1 = -3.048846467e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = 4.440892099e-22 ppdiblc1 = -5.551115123e-29
+ pdiblc2 = -8.673906562e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 1.301042607e-23 ppdiblc2 = -1.084202172e-31
+ pdiblcb = -8.553970445e-02 lpdiblcb = -4.630533311e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076329e+07 lpscbe1 = 1.888714223e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729690e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380752e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373076e+03 lat = 9.625574770e-3
+ ute = -1.301136473e+00 lute = -4.669823644e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393852e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873018e-25 wub1 = 6.162975822e-39 pub1 = -1.540743956e-45
+ uc1 = -1.418079324e-10 luc1 = 7.536563684e-17 wuc1 = 2.067951531e-31 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.115 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.910376278e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456612608e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016978168e-18
+ cit = 0.0
+ voff = {-9.930380979e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149569577e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935962584e-16
+ ags = 1.250000000e+00 lags = 6.286171583e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-08 wketa = -8.881784197e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026379313e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347644218e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990585640e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.630233765e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009865197e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190619704e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.116 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {8.061145465e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.325626486e-08 wvth0 = -8.114210699e-08 pvth0 = 1.548077803e-14
+ k1 = 0.90707349
+ k2 = -1.872942668e-01 lk2 = 8.178558149e-09 wk2 = 4.302656511e-08 pk2 = -8.208866250e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.584992040e-01 ldsub = 2.495405448e-11 wdsub = 6.961098779e-11 pdsub = -1.328080192e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079725281e-19
+ cit = 0.0
+ voff = {-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.724220849e-17
+ nfactor = 1.334758330e+01 lnfactor = -2.179648517e-06 wnfactor = -6.044194464e-06 pnfactor = 1.153147685e-12
+ eta0 = 1.826779867e-02 leta0 = -3.485240187e-09 weta0 = -9.717226783e-09 peta0 = 1.853910829e-15
+ etab = -0.043998
+ u0 = -8.465704720e-02 lu0 = 2.109378145e-08 wu0 = 6.413598440e-08 pu0 = -1.223624792e-14
+ ua = -3.087979294e-09 lua = 3.806657188e-16 wua = 1.045373434e-15 pua = -1.994426159e-22
+ ub = 2.653968253e-17 lub = -4.791789839e-24 wub = -1.324030475e-23 pub = 2.526064782e-30
+ uc = 3.550112941e-10 luc = -5.303989961e-17 wuc = -1.479585772e-16 puc = 2.822842511e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.914970573e+05 lvsat = 1.490802965e-01 wvsat = 2.094686876e-01 pvsat = -3.996369303e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.325212843e-05 lb0 = 2.525359119e-12 wb0 = 6.996719441e-12 pb0 = -1.334876115e-18
+ b1 = 2.663317764e-06 lb1 = -5.060953252e-13 wb1 = -1.380737492e-12 pb1 = 2.634253832e-19
+ keta = -2.700000009e-02 lketa = 1.434297126e-17
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.564208446e-01 lpclm = 1.022010321e-07 wpclm = 2.743800111e-07 ppclm = -5.234786480e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.150327289e-24
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968377e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.983091288e-01 lkt1 = 5.088104192e-08 wkt1 = 1.399896776e-07 pkt1 = -2.670807063e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.578778028e-11
+ ute = 3.963587508e-01 lute = -3.266482377e-07 wute = -9.018427563e-07 pute = 1.720589721e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.117 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.118 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.549167264e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016575863e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = 7.629394531e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.119 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.031067740e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-07 pk2 = 2.220446049e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179965467e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647567e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = 4.440892099e-22 ppclm = -2.664535259e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267871e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15 wua1 = 3.308722450e-30
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16 wuc1 = -5.169878828e-32 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.120 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.427426575e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-06 wdsub = -1.776356839e-21
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.375696972e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14 wb0 = -1.058791184e-28
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14 pb1 = 2.646977960e-35
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.121 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.911229542e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.358925766e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159063e-03 leta0 = 4.128463499e-09 weta0 = -1.734723476e-24
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -3.295974604e-23 petab = 4.163336342e-29
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24 pub = -1.540743956e-45
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-06 pags = -1.776356839e-27
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 wb0 = 5.293955920e-29 pb0 = 5.293955920e-35
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = 2.775557562e-23 pketa = -2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 7.411538288e-28 palpha0 = 4.976318565e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -1.240770919e-30 pua1 = -8.271806126e-37
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 pub1 = -7.703719778e-46
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.122 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.821975320e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.303523806e-08 wvth0 = 3.447097530e-08 pvth0 = -3.484277924e-14
+ k1 = 6.351021960e-01 lk1 = -8.178610772e-08 wk1 = -3.526778869e-16 pk1 = 3.564819551e-22
+ k2 = -9.819090370e-02 lk2 = 5.532097549e-08 wk2 = 8.890189169e-09 pk2 = -8.986078750e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076448e-01 ldsub = 5.194667313e-08 wdsub = -1.040207920e-16 pdsub = 1.051430054e-22
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.255026654e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.262473516e-09 wvoff = -4.291291766e-16 pvoff = 4.337576964e-22
+ nfactor = 1.616966924e+00 lnfactor = 6.097217582e-07 wnfactor = -4.169514511e-15 pnfactor = 4.214484761e-21
+ eta0 = -4.954531764e-01 leta0 = 5.033556864e-07 weta0 = 2.379968514e-16 peta0 = -2.405640999e-22
+ etab = -1.699316551e-01 letab = 8.647946918e-08 wetab = 4.781841589e-17 petab = -4.833422551e-23
+ u0 = -2.210078630e-03 lu0 = 2.447848620e-08 wu0 = 1.361929054e-08 pu0 = -1.376618821e-14
+ ua = -6.439294864e-10 lua = -4.848815377e-16 wua = 2.370166855e-21 pua = -2.395731474e-27
+ ub = 1.111498246e-18 lub = 2.659901090e-25 wub = 2.370352916e-30 pub = -2.395919541e-36
+ uc = 2.628890927e-11 luc = 1.340715722e-17 wuc = -5.360678376e-26 puc = 5.418487962e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.914931349e+06 lvsat = 3.030687524e+00 wvsat = 1.323176037e+00 pvsat = -1.337447814e-6
+ a0 = 1.011417803e+00 la0 = 1.906162443e-07 wa0 = 2.592706494e-15 pa0 = -2.620669903e-21
+ ags = 2.367344351e+00 lags = -1.129396027e-06 wags = 1.145646067e-14 pags = -1.158003116e-20
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907885e-08 lb0 = -1.871983642e-14 wb0 = -2.718684593e-23 pb0 = 2.748010462e-29
+ b1 = 6.204608816e-08 lb1 = -3.169227335e-14 wb1 = -1.572521961e-22 pb1 = 1.589483266e-28
+ keta = -1.194413453e-01 lketa = 5.737558669e-08 wketa = 3.952973504e-16 pketa = -3.995610509e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898536e+00 lpclm = -4.321701819e-07 wpclm = -3.028485906e-15 ppclm = 3.061151332e-21
+ pdiblc1 = 6.826367982e-01 lpdiblc1 = -3.318091416e-07 wpdiblc1 = 5.676632497e-16 ppdiblc1 = -5.737854636e-22
+ pdiblc2 = 9.443109138e-03 lpdiblc2 = -4.799688249e-09 wpdiblc2 = -1.368019587e-17 ppdiblc2 = 1.382775838e-23
+ pdiblcb = 9.625889866e-02 lpdiblcb = -9.749071449e-08 wpdiblcb = 1.099100186e-16 ppdiblcb = -1.110955247e-22
+ drout = 8.376749873e-01 ldrout = 8.291329245e-08 wdrout = -3.815046057e-16 pdrout = 3.856222008e-22
+ pscbe1 = 1.037253089e+09 lpscbe1 = -3.066279363e+02 wpscbe1 = 4.392906189e-06 ppscbe1 = -4.440286636e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946629e-06 lalpha0 = -1.672796883e-12 walpha0 = 5.156357112e-21 palpha0 = -5.211976684e-27
+ alpha1 = 0.85
+ beta0 = 1.689804916e+01 lbeta0 = 5.720551851e-07 wbeta0 = -2.295894319e-14 pbeta0 = 2.320655312e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718610e-01 lkt1 = -4.432457352e-09 wkt1 = 3.684341721e-17 pkt1 = -3.724087705e-23
+ kt2 = -1.732617330e-02 lkt2 = -9.905380060e-09 wkt2 = 6.005085318e-18 pkt2 = -6.069811320e-24
+ at = 1.158432499e+05 lat = -5.372855215e-02 wat = 4.562644754e-10 pat = -4.611859331e-16
+ ute = -8.338566420e-01 lute = -2.433498205e-07 wute = -9.430962677e-16 pute = 9.532676870e-22
+ ua1 = 1.741162740e-09 lua1 = -4.645563762e-16 wua1 = 1.953780755e-24 pua1 = -1.974854008e-30
+ ub1 = -7.096737815e-19 lub1 = 3.973648573e-26 wub1 = 4.286565388e-34 pub1 = -4.332787707e-40
+ uc1 = 7.705161076e-11 luc1 = -3.642475380e-17 wuc1 = -4.747582446e-26 puc1 = 4.798784926e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.123 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {7.776929907e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.789970531e-08 wvth0 = -6.894195061e-08 pvth0 = 1.797909553e-14
+ k1 = 2.425254185e-02 lk1 = 2.302273437e-07 wk1 = 7.053557738e-16 pk1 = -1.839470798e-22
+ k2 = 1.741672963e-01 lk2 = -8.379578003e-08 wk2 = -1.778037834e-08 pk2 = 4.636873745e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850176e-01 ldsub = 7.902988878e-08 wdsub = 2.080424721e-16 pdsub = -5.425460081e-23
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
+ voff = {-1.072895709e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.856546724e-08 wvoff = 8.582583533e-16 pvoff = -2.238217389e-22
+ nfactor = 4.181852111e+00 lnfactor = -7.003856872e-07 wnfactor = 8.339029023e-15 pnfactor = -2.174701308e-21
+ eta0 = 1.000416473e+00 leta0 = -2.607135883e-07 weta0 = -4.759943550e-16 peta0 = 1.241322600e-22
+ etab = 4.461928492e-02 letab = -2.311014727e-08 wetab = -9.563704863e-17 petab = 2.494078381e-23
+ u0 = 7.223690378e-02 lu0 = -1.354799016e-08 wu0 = -2.723858107e-08 pu0 = 7.103440604e-15
+ ua = -2.102021197e-09 lua = 2.598912947e-16 wua = -4.740333710e-21 pua = 1.236212667e-27
+ ub = 2.286040547e-18 lub = -3.339496549e-25 wub = -4.740705826e-30 pub = 1.236309710e-36
+ uc = 1.078724744e-11 luc = 2.132518905e-17 wuc = 1.072133607e-25 puc = -2.795979038e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.882720731e+06 lvsat = -1.463029992e+00 wvsat = -2.646352074e+00 pvsat = 6.901315721e-7
+ a0 = 1.264221194e+00 la0 = 6.148781164e-08 wa0 = -5.185412988e-15 pa0 = 1.352281842e-21
+ ags = -9.846887014e-01 lags = 5.827755276e-07 wags = -2.291292400e-14 pags = 5.975369533e-21
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.152151564e-16 lb0 = 3.004649978e-23 wb0 = 5.437371919e-23 pb0 = -1.417990473e-29
+ b1 = -6.664189737e-16 lb1 = 1.737927385e-22 wb1 = 3.145044391e-22 pb1 = -8.201835465e-29
+ keta = 7.220181600e-02 lketa = -4.051305711e-08 wketa = -7.905947008e-16 pketa = 2.061760276e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500137e-01 lpclm = -1.136192480e-07 wpclm = 6.056973589e-15 ppclm = -1.579573805e-21
+ pdiblc1 = -3.048846444e-01 lpdiblc1 = 1.726029860e-07 wpdiblc1 = -1.135325833e-15 ppdiblc1 = 2.960770240e-22
+ pdiblc2 = -8.673906618e-03 lpdiblc2 = 4.454229761e-09 wpdiblc2 = 2.736040409e-17 ppdiblc2 = -7.135207789e-24
+ pdiblcb = -8.553970401e-02 lpdiblcb = -4.630533427e-09 wpdiblcb = -2.198201621e-16 ppdiblcb = 5.732603281e-23
+ drout = 1.518101609e+00 ldrout = -2.646391000e-07 wdrout = 7.630127641e-16 pdrout = -1.989830523e-22
+ pscbe1 = 6.718078115e+07 lpscbe1 = 1.888714176e+02 wpscbe1 = -8.785812378e-06 ppscbe1 = 2.291216850e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729711e-06 lalpha0 = -2.066502091e-12 walpha0 = -1.031272778e-20 palpha0 = 2.689410923e-27
+ alpha1 = 0.85
+ beta0 = 2.187554641e+01 lbeta0 = -1.970380727e-06 wbeta0 = 4.591782954e-14 pbeta0 = -1.197473409e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774103e-01 lkt1 = 2.024134099e-08 wkt1 = -7.368683441e-17 pkt1 = 1.921640624e-23
+ kt2 = -4.489649531e-02 lkt2 = 4.177154438e-09 wkt2 = -1.201017064e-17 pkt2 = 3.132077930e-24
+ at = -8.189371221e+03 lat = 9.625574286e-03 wat = -9.125292418e-10 pat = 2.379748476e-16
+ ute = -1.301136477e+00 lute = -4.669822644e-09 wute = 1.886192535e-15 pute = -4.918909724e-22
+ ua1 = 1.724096906e-09 lua1 = -4.558393872e-16 wua1 = -3.907558200e-24 pua1 = 1.019036057e-30
+ ub1 = -2.029308258e-18 lub1 = 7.137873014e-25 wub1 = -8.573099962e-34 pub1 = 2.235750443e-40
+ uc1 = -1.418079326e-10 luc1 = 7.536563689e-17 wuc1 = 9.495149383e-26 puc1 = -2.476198768e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.124 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.910376278e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456790244e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
+ voff = {-9.930380979e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149680599e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935927057e-16
+ ags = 1.250000000e+00 lags = 6.285816312e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026201677e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347671974e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990363595e-18
+ drout = 5.033266586e-01 ldrout = 2.662101650e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.630043030e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009865197e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.191033295e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.125 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {9.627035343e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.313125148e-08 wvth0 = -1.581732409e-07 pvth0 = 3.017723995e-14
+ k1 = 0.90707349
+ k2 = -4.976247873e-01 lk2 = 6.738527684e-08 wk2 = 1.956880787e-07 pk2 = -3.733454579e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585002188e-01 ldsub = 2.476043415e-11 wdsub = 6.911174762e-11 pdsub = -1.318555388e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079655892e-19
+ cit = 0.0
+ voff = {-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.724309667e-17
+ nfactor = 1.334758404e+01 lnfactor = -2.179648659e-06 wnfactor = -6.044194829e-06 pnfactor = 1.153147755e-12
+ eta0 = 1.826779849e-02 leta0 = -3.485240153e-09 weta0 = -9.717226695e-09 peta0 = 1.853910812e-15
+ etab = -0.043998
+ u0 = 4.637763925e-01 lu0 = -8.353964079e-08 wu0 = -2.056559745e-07 pu0 = 3.923628075e-14
+ ua = -3.087976251e-09 lua = 3.806651381e-16 wua = 1.045371936e-15 pua = -1.994423302e-22
+ ub = 2.653990193e-17 lub = -4.791831698e-24 wub = -1.324041268e-23 pub = 2.526085373e-30
+ uc = 3.528542115e-10 luc = -5.262835845e-17 wuc = -1.468974392e-16 puc = 2.802597484e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.016421737e+06 lvsat = 1.203158576e+00 wvsat = 2.927355935e+00 pvsat = -5.584985294e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.325201989e-05 lb0 = 2.525338411e-12 wb0 = 6.996666048e-12 pb0 = -1.334865929e-18
+ b1 = 2.663305599e-06 lb1 = -5.060930044e-13 wb1 = -1.380731508e-12 pb1 = 2.634242415e-19
+ keta = -2.700000009e-02 lketa = 1.434308228e-17
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.564201645e-01 lpclm = 1.022009023e-07 wpclm = 2.743796765e-07 ppclm = -5.234780096e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.150539047e-24
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968377e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.983091390e-01 lkt1 = 5.088104389e-08 wkt1 = 1.399896827e-07 pkt1 = -2.670807160e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.578824595e-11
+ ute = 3.832108188e-01 lute = -3.241397963e-07 wute = -8.953748678e-07 pute = 1.708249895e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.126 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.127 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.549167264e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.252285745e-7
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016575863e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-07 wa0 = 1.776356839e-21
+ ags = 3.207608585e-01 lags = 4.826429794e-07 wags = -4.440892099e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.128 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.031067740e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-07 pk2 = -1.110223025e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179965467e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647566e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-08 pketa = -5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 ppclm = 3.108624469e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267871e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.129 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.427426575e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.375696972e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.130 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.911229542e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.358925766e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159063e-03 leta0 = 4.128463499e-09 weta0 = 8.673617380e-25
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -4.336808690e-24 petab = -6.938893904e-30
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15 pua = 8.271806126e-37
+ ub = -2.930959084e-19 lub = 1.685734216e-24
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-06 pags = 8.881784197e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 wb0 = 5.293955920e-29 pb0 = 5.293955920e-35
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = -1.387778781e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 2.805796638e-27 palpha0 = -1.799945013e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = 4.135903063e-31 pua1 = -1.654361225e-36
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 wub1 = -3.851859889e-40 pub1 = -3.851859889e-46
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.131 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.552397824e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.920515398e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610696e-8
+ k2 = -7.935304322e-02 lk2 = 3.627992986e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667335e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.255026664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.262472597e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217672e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -7.632783294e-23 peta0 = 1.214306433e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.664850807e-02 lu0 = -4.691369216e-9
+ ua = -6.439244642e-10 lua = -4.848866142e-16
+ ub = 1.111503269e-18 lub = 2.659850321e-25
+ uc = 2.628890915e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.111883581e+05 lvsat = 1.967033607e-01 pvsat = 1.164153218e-22
+ a0 = 1.011417809e+00 la0 = 1.906162387e-7
+ ags = 2.367344375e+00 lags = -1.129396051e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608782e-08 lb1 = -3.169227302e-14
+ keta = -1.194413445e-01 lketa = 5.737558585e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701755e-7
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109109e-03 lpdiblc2 = -4.799688220e-9
+ pdiblcb = 9.625889889e-02 lpdiblcb = -9.749071473e-08 wpdiblcb = -1.908195824e-23 ppdiblcb = -2.146720302e-29
+ drout = 8.376749865e-01 ldrout = 8.291329327e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279457e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552343e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457430e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380073e-9
+ at = 1.158432509e+05 lat = -5.372855313e-2
+ ute = -8.338566440e-01 lute = -2.433498184e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563804e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648481e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475369e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.132 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.316084900e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.980291269e-8
+ k1 = 2.425254334e-02 lk1 = 2.302273434e-7
+ k2 = 1.364915753e-01 lk2 = -7.397047947e-08 wk2 = 2.775557562e-23 pk2 = 5.204170428e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988866e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
+ voff = {-1.072895691e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.856546771e-8
+ nfactor = 4.181852129e+00 lnfactor = -7.003856918e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928472e-02 letab = -2.311014721e-08 wetab = -6.938893904e-24 petab = 1.214306433e-29
+ u0 = 1.451973038e-02 lu0 = 1.503840623e-9
+ ua = -2.102031242e-09 lua = 2.598939142e-16
+ ub = 2.286030502e-18 lub = -3.339470352e-25
+ uc = 1.078724767e-11 luc = 2.132518899e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.752347497e+05 lvsat = -6.761528150e-4
+ a0 = 1.264221183e+00 la0 = 6.148781451e-8
+ ags = -9.846887499e-01 lags = 5.827755403e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.220181432e-02 lketa = -4.051305667e-08 wketa = 1.387778781e-23 pketa = -1.734723476e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500265e-01 lpclm = -1.136192514e-7
+ pdiblc1 = -3.048846468e-01 lpdiblc1 = 1.726029866e-07 ppdiblc1 = 6.938893904e-29
+ pdiblc2 = -8.673906560e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 3.252606517e-25 ppdiblc2 = -3.523657061e-31
+ pdiblcb = -8.553970447e-02 lpdiblcb = -4.630533306e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076254e+07 lpscbe1 = 1.888714225e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729689e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380753e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-08 wkt1 = 4.440892099e-22
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373154e+03 lat = 9.625574790e-3
+ ute = -1.301136473e+00 lute = -4.669823687e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393851e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873019e-25
+ uc1 = -1.418079323e-10 luc1 = 7.536563684e-17 wuc1 = 5.169878828e-32 puc1 = 2.261821987e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.133 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.910376278e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456701426e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
+ voff = {-9.930380979e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149680599e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935962584e-16
+ ags = 1.250000000e+00 lags = 6.285993948e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026201677e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347658096e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990363595e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.630043030e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009864680e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190826499e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.134 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {1.640247921e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.023972348e-07 wvth0 = -4.779281183e-07 pvth0 = 9.118199398e-14
+ k1 = 0.90707349
+ k2 = -3.443785481e-01 lk2 = 3.814803985e-08 wk2 = 1.233662746e-07 pk2 = -2.353655806e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585021073e-01 ldsub = 2.440014616e-11 wdsub = 6.822053216e-11 pdsub = -1.301552245e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079517114e-19
+ cit = 0.0
+ voff = {-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.724309667e-17
+ nfactor = 1.334758347e+01 lnfactor = -2.179648551e-06 wnfactor = -6.044194562e-06 pnfactor = 1.153147704e-12
+ eta0 = 1.826777218e-02 leta0 = -3.485235134e-09 weta0 = -9.717214281e-09 peta0 = 1.853908444e-15
+ etab = -0.043998
+ u0 = 2.066270621e-01 lu0 = -3.447914862e-08 wu0 = -8.429897664e-08 pu0 = 1.608306456e-14
+ ua = -3.087977982e-09 lua = 3.806654685e-16 wua = 1.045372754e-15 pua = -1.994424862e-22
+ ub = 2.653983749e-17 lub = -4.791819404e-24 wub = -1.324038227e-23 pub = 2.526079571e-30
+ uc = 3.488330108e-10 luc = -5.186116966e-17 wuc = -1.449997060e-16 puc = 2.766391390e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.128720330e+06 lvsat = 8.430115758e-01 wvsat = 2.036489235e+00 pvsat = -3.885336351e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.325205743e-05 lb0 = 2.525345573e-12 wb0 = 6.996683763e-12 pb0 = -1.334869308e-18
+ b1 = 2.663308614e-06 lb1 = -5.060935796e-13 wb1 = -1.380732931e-12 pb1 = 2.634245130e-19
+ keta = -2.700000009e-02 lketa = 1.434302677e-17
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.564203852e-01 lpclm = 1.022009444e-07 wpclm = 2.743797807e-07 ppclm = -5.234782084e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -3.150539047e-24
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968377e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.983091505e-01 lkt1 = 5.088104606e-08 wkt1 = 1.399896881e-07 pkt1 = -2.670807262e-14
+ kt2 = -0.028878939
+ at = 5.372048690e+04 lat = 1.578801312e-11
+ ute = 3.587006802e-01 lute = -3.194636050e-07 wute = -8.838077490e-07 pute = 1.686181452e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.135 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.136 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.549167264e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.252285745e-07 wvth0 = 1.776356839e-21
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016575863e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-07 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = 7.629394531e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16 puc1 = -1.654361225e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.137 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.031067740e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179965467e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647567e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = -4.440892099e-22 ppclm = -7.105427358e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-08 ppdiblc2 = -2.775557562e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267872e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16 puc1 = 8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.138 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.427426575e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.375696972e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14 wb0 = 2.117582368e-28
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-06 wpclm = -3.552713679e-21
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.139 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.911229542e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.358925766e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-6
+ eta0 = -1.553159063e-03 leta0 = 4.128463499e-09 peta0 = 3.469446952e-30
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = -1.734723476e-23 petab = 1.075528555e-28
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24 pub = -3.081487911e-45
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 wb0 = -1.058791184e-28 pb0 = -1.058791184e-34
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = -1.110223025e-22 pketa = -1.665334537e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = 6.564505341e-27 palpha0 = -4.235164736e-34
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -1.654361225e-30
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 wub1 = -7.703719778e-40 pub1 = 2.311115933e-45
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.140 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.552397824e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.920515398e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610696e-8
+ k2 = -7.935304322e-02 lk2 = 3.627992986e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667335e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.255026664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.262472597e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217672e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 2.498001805e-22 peta0 = -1.387778781e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.664850807e-02 lu0 = -4.691369216e-9
+ ua = -6.439244642e-10 lua = -4.848866142e-16
+ ub = 1.111503269e-18 lub = 2.659850321e-25
+ uc = 2.628890915e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.111883581e+05 lvsat = 1.967033607e-1
+ a0 = 1.011417809e+00 la0 = 1.906162387e-7
+ ags = 2.367344375e+00 lags = -1.129396051e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608782e-08 lb1 = -3.169227302e-14
+ keta = -1.194413445e-01 lketa = 5.737558585e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701755e-7
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109109e-03 lpdiblc2 = -4.799688220e-9
+ pdiblcb = 9.625889889e-02 lpdiblcb = -9.749071473e-08 wpdiblcb = 1.023486851e-22 ppdiblcb = 6.028164079e-29
+ drout = 8.376749865e-01 ldrout = 8.291329327e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279457e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552343e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457430e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380073e-9
+ at = 1.158432509e+05 lat = -5.372855313e-2
+ ute = -8.338566440e-01 lute = -2.433498184e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563804e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648481e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475369e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.141 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.316084900e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.980291269e-8
+ k1 = 2.425254334e-02 lk1 = 2.302273434e-7
+ k2 = 1.364915753e-01 lk2 = -7.397047947e-08 wk2 = -1.665334537e-22 pk2 = -9.714451465e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988866e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
+ voff = {-1.072895691e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.856546771e-8
+ nfactor = 4.181852129e+00 lnfactor = -7.003856918e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928472e-02 letab = -2.311014721e-08 wetab = 4.857225733e-23 petab = -1.387778781e-29
+ u0 = 1.451973038e-02 lu0 = 1.503840623e-9
+ ua = -2.102031242e-09 lua = 2.598939142e-16
+ ub = 2.286030502e-18 lub = -3.339470352e-25
+ uc = 1.078724767e-11 luc = 2.132518899e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.752347497e+05 lvsat = -6.761528150e-4
+ a0 = 1.264221183e+00 la0 = 6.148781451e-8
+ ags = -9.846887499e-01 lags = 5.827755403e-07 wags = 1.776356839e-21 pags = -4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.220181432e-02 lketa = -4.051305667e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500265e-01 lpclm = -1.136192514e-7
+ pdiblc1 = -3.048846468e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = 4.440892099e-22 ppdiblc1 = -1.110223025e-28
+ pdiblc2 = -8.673906560e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = -4.119968255e-24 ppdiblc2 = -5.854691731e-30
+ pdiblcb = -8.553970447e-02 lpdiblcb = -4.630533306e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076254e+07 lpscbe1 = 1.888714225e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729689e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380753e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373154e+03 lat = 9.625574790e-03 pat = 1.455191523e-23
+ ute = -1.301136473e+00 lute = -4.669823687e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393851e-16 wua1 = -6.617444900e-30
+ ub1 = -2.029308260e-18 lub1 = 7.137873019e-25 pub1 = -7.703719778e-46
+ uc1 = -1.418079323e-10 luc1 = 7.536563684e-17 wuc1 = -2.584939414e-32 puc1 = 6.462348536e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.142 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.910376278e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610801044e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456790244e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016992046e-18
+ cit = 0.0
+ voff = {-9.930380979e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.150013666e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935820476e-16
+ ags = 1.250000000e+00 lags = 6.286882126e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026379313e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347644218e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990585640e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629852295e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009866231e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190619704e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.143 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {-2.712151192e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.279795823e-07 wvth0 = 1.445536326e-06 pvth0 = -2.757880936e-13
+ k1 = 0.90707349
+ k2 = 2.080083157e-01 lk2 = -6.723964035e-08 wk2 = -1.207511569e-07 pk2 = 2.303763022e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.687830613e+00 ldsub = -4.253002681e-07 wdsub = -9.851433845e-07 pdsub = 1.879515657e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079586503e-19
+ cit = 0.0
+ voff = {-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.724220849e-17
+ nfactor = -3.997886150e+00 lnfactor = 1.129624217e-06 wnfactor = 1.621323520e-06 pnfactor = -3.093258290e-13
+ eta0 = -1.264688194e-02 leta0 = 2.412848068e-09 weta0 = 3.944960646e-09 peta0 = -7.526432618e-16
+ etab = -0.043998
+ u0 = 4.427431561e-01 lu0 = -7.952679374e-08 wu0 = -1.886462343e-07 pu0 = 3.599106046e-14
+ ua = -1.023251079e-09 lua = -1.325551842e-17 wua = 1.329038639e-16 pua = -2.535619658e-23
+ ub = -4.555577596e-18 lub = 1.140750460e-24 wub = 5.016767147e-25 pub = -9.571289368e-32
+ uc = -2.391896018e-10 luc = 6.032531251e-17 wuc = 1.148663033e-16 puc = -2.191488254e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.313909858e+06 lvsat = -9.585100672e-01 wvsat = -2.136511210e+00 pvsat = 4.076164276e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.404797633e-06 lb0 = -6.525491778e-13 wb0 = -3.645135095e-13 pb0 = 6.954407442e-20
+ b1 = 2.644971507e-06 lb1 = -5.025951163e-13 wb1 = -1.372629177e-12 pb1 = 2.618784301e-19
+ keta = -8.680480736e-01 lketa = 1.604601978e-07 wketa = 3.716860572e-07 pketa = -7.091249611e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.238634796e-02 lpclm = 3.183778305e-08 wpclm = 1.113922835e-07 ppclm = -2.125208819e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.999997308e-08 lalpha0 = 5.135634875e-21 walpha0 = 1.190335528e-20 palpha0 = -2.270993587e-27
+ alpha1 = 0.85
+ beta0 = 1.393352495e+01 lbeta0 = -1.342963468e-08 wbeta0 = 1.137225354e-13 pbeta0 = -2.169667823e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.815416568e-01 lkt1 = -9.553756987e-09 wkt1 = -3.972203899e-15 pkt1 = 7.578409011e-22
+ kt2 = -0.028878939
+ at = 5.372048980e+04 lat = -5.378732458e-10 wat = -1.282487996e-09 pat = 2.446807921e-16
+ ute = -1.155115866e+00 lute = -3.064860140e-08 wute = -2.148037751e-07 pute = 4.098155304e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.144 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.145 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.549167264e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.252285745e-07 wvth0 = -8.881784197e-22
+ k1 = 6.125245790e-01 lk1 = -8.908173397e-7
+ k2 = -4.542695903e-02 lk2 = 2.699597714e-07 pk2 = 4.440892099e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016575863e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.324764808e-7
+ nfactor = 4.357652976e+00 lnfactor = -8.713756309e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952409390e-02 lu0 = 4.963087355e-8
+ ua = -1.237271306e-09 lua = 3.764549248e-15
+ ub = 1.292509458e-18 lub = -8.836654604e-25
+ uc = 6.336963784e-11 luc = -2.968127417e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.391038290e+00 la0 = -5.690725414e-7
+ ags = 3.207608585e-01 lags = 4.826429794e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.182065634e-08 lb0 = -4.969365854e-14
+ b1 = 1.716224571e-08 lb1 = -9.579654950e-14
+ keta = -2.652182624e-03 lketa = -3.790878070e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.827620000e-03 lpclm = 5.343404145e-07 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.498814613e-04 lpdiblc2 = 8.213347045e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.540394762e+07 lpscbe1 = 6.011319109e+03 ppscbe1 = 3.814697266e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832023882e-01 lkt1 = -6.358650932e-8
+ kt2 = -3.549038051e-02 lkt2 = 1.195134091e-7
+ at = 1.983647925e+05 lat = -4.675478627e-1
+ ute = -1.015465445e+00 lute = -1.999769001e-6
+ ua1 = 1.029476770e-09 lua1 = 1.831451771e-15
+ ub1 = -3.818573919e-19 lub1 = -3.754275752e-24
+ uc1 = 6.946434833e-11 luc1 = -7.133042041e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.146 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.031067740e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.391884164e-7
+ k1 = 4.363871732e-01 lk1 = 5.201817251e-7
+ k2 = 2.091918684e-02 lk2 = -2.615250051e-07 pk2 = -1.110223025e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179965467e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.588565194e-9
+ nfactor = 3.994589269e+00 lnfactor = -5.805330654e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.371290349e-02 lu0 = 1.607521627e-8
+ ua = -9.745240495e-10 lua = 1.659737204e-15
+ ub = 1.352036733e-18 lub = -1.360525724e-24
+ uc = 9.453647566e-12 luc = 1.350967184e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.410242685e+00 la0 = -7.229148376e-7
+ ags = 3.607956386e-01 lags = 1.619329236e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.293006201e-09 lb0 = -1.340284109e-13
+ b1 = 6.090685054e-09 lb1 = -7.104646376e-15
+ keta = -1.755174251e-02 lketa = 8.144840504e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.011084057e-01 lpclm = 6.072042855e-06 wpclm = 2.220446049e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.671405040e-03 lpdiblc2 = 2.600759785e-08 ppdiblc2 = -1.387778781e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.386978466e+08 lpscbe1 = 2.908024536e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862267871e-01 lkt1 = -3.935869671e-8
+ kt2 = -9.701244670e-03 lkt2 = -8.707783927e-8
+ at = 140000.0
+ ute = -1.230707510e+00 lute = -2.755108770e-7
+ ua1 = 1.518149337e-09 lua1 = -2.083199590e-15
+ ub1 = -1.029000004e-18 lub1 = 1.429845225e-24
+ uc1 = -7.165275628e-11 luc1 = 4.171547218e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.147 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.427426575e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.978263048e-8
+ k1 = 5.590290829e-01 lk1 = 2.829127054e-8
+ k2 = -4.522950576e-02 lk2 = 3.783245109e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.616179000e-01 ldsub = -1.209724851e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.375696972e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.691515281e-8
+ nfactor = 1.874008369e+00 lnfactor = 2.699865535e-6
+ eta0 = 1.599287435e-01 leta0 = -3.205770854e-7
+ etab = -1.398748135e-01 letab = 2.802529237e-7
+ u0 = 2.954679423e-02 lu0 = -7.323271004e-9
+ ua = -7.063921832e-10 lua = 5.843176682e-16
+ ub = 1.482911605e-18 lub = -1.885436828e-24
+ uc = 3.544272737e-11 luc = 3.086008094e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.617277384e+00 la0 = -1.553286708e-6
+ ags = 3.254840150e-01 lags = 3.035602892e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.052382650e-08 lb0 = 6.342587392e-14
+ b1 = -6.790996425e-09 lb1 = 4.456102136e-14
+ keta = 4.786864729e-04 lketa = 9.132212898e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.121656622e+00 lpclm = -1.238677599e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.433178216e-03 lpdiblc2 = 9.544992792e-9
+ pdiblcb = -3.756741250e-02 lpdiblcb = 5.040520211e-8
+ drout = 0.56
+ pscbe1 = 6.219270175e+08 lpscbe1 = 3.580666602e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.580562525e-01 lkt1 = -1.523446829e-7
+ kt2 = -1.446881568e-02 lkt2 = -6.795613219e-8
+ at = 1.707951876e+05 lat = -1.235129073e-1
+ ute = -8.660756170e-01 lute = -1.737971369e-6
+ ua1 = 2.160350910e-09 lua1 = -4.658932669e-15
+ ub1 = -1.500370758e-18 lub1 = 3.320412446e-24 pub1 = 3.081487911e-45
+ uc1 = 7.997501133e-12 luc1 = 9.769458448e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.148 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.911229542e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.401354624e-8
+ k1 = 5.922128235e-01 lk1 = -3.843413038e-8
+ k2 = -4.323459656e-02 lk2 = -2.280903676e-10
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.358925766e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.184367932e-8
+ nfactor = 4.223966039e+00 lnfactor = -2.025396449e-06 wnfactor = 7.105427358e-21
+ eta0 = -1.553159062e-03 leta0 = 4.128463499e-9
+ etab = 8.427967575e-02 letab = -1.704737851e-07 wetab = 1.561251128e-23 petab = 1.110223025e-28
+ u0 = 2.984443951e-02 lu0 = -7.921771979e-9
+ ua = 2.996706033e-10 lua = -1.438659298e-15
+ ub = -2.930959084e-19 lub = 1.685734216e-24
+ uc = 6.214820228e-11 luc = -2.283891413e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.654715502e+04 lvsat = 6.942932338e-3
+ a0 = 4.857688128e-01 la0 = 7.219348848e-7
+ ags = -3.054435103e-01 lags = 1.572220524e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.649126846e-08 lb0 = 7.542512268e-14 wb0 = -5.293955920e-29
+ b1 = -1.172630920e-10 lb1 = 3.114157180e-14
+ keta = 7.344880195e-02 lketa = -1.375950737e-07 wketa = -2.775557562e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.370063458e-01 lpclm = 7.412433910e-7
+ pdiblc1 = 4.260159629e-01 lpdiblc1 = -7.242039391e-8
+ pdiblc2 = 9.692319220e-03 lpdiblc2 = -5.051586311e-9
+ pdiblcb = -2.494125765e-02 lpdiblcb = 2.501670671e-8
+ drout = 1.964167178e-01 ldrout = 7.310881736e-7
+ pscbe1 = 8.668158353e+08 lpscbe1 = -1.343523463e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.519215140e-06 lalpha0 = 1.115828411e-11 walpha0 = -5.293955920e-28 palpha0 = -5.717472394e-33
+ alpha1 = 0.85
+ beta0 = 1.021712726e+01 lbeta0 = 7.325037513e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.936211119e-01 lkt1 = 1.202472386e-7
+ kt2 = -6.963139074e-02 lkt2 = 4.296400146e-8
+ at = 1.565554817e+05 lat = -9.487990606e-2
+ ute = -2.393263654e+00 lute = 1.332876956e-6
+ ua1 = -1.610315848e-09 lua1 = 2.923071260e-15 wua1 = -4.135903063e-31 pua1 = 4.135903063e-37
+ ub1 = 9.810797682e-19 lub1 = -1.669253532e-24 wub1 = -3.851859889e-40 pub1 = -1.540743956e-45
+ uc1 = 7.231791215e-11 luc1 = -3.163999752e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.149 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.552397824e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.920515398e-8
+ k1 = 6.351021953e-01 lk1 = -8.178610696e-8
+ k2 = -7.935304322e-02 lk2 = 3.627992986e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.086076446e-01 ldsub = 5.194667335e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.255026664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.262472597e-9
+ nfactor = 1.616966915e+00 lnfactor = 6.097217672e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -2.081668171e-22 peta0 = 2.810252031e-28
+ etab = -1.699316550e-01 letab = 8.647946908e-8
+ u0 = 2.664850807e-02 lu0 = -4.691369216e-9
+ ua = -6.439244642e-10 lua = -4.848866142e-16
+ ub = 1.111503269e-18 lub = 2.659850321e-25
+ uc = 2.628890915e-11 luc = 1.340715733e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.111883581e+05 lvsat = 1.967033607e-01 pvsat = -1.164153218e-22
+ a0 = 1.011417809e+00 la0 = 1.906162387e-7
+ ags = 2.367344375e+00 lags = -1.129396051e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.664907879e-08 lb0 = -1.871983636e-14
+ b1 = 6.204608782e-08 lb1 = -3.169227302e-14
+ keta = -1.194413445e-01 lketa = 5.737558585e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.297898529e+00 lpclm = -4.321701755e-7
+ pdiblc1 = 6.826367994e-01 lpdiblc1 = -3.318091428e-7
+ pdiblc2 = 9.443109109e-03 lpdiblc2 = -4.799688220e-9
+ pdiblcb = 9.625889889e-02 lpdiblcb = -9.749071473e-08 wpdiblcb = 4.336808690e-24 ppdiblcb = 2.016616041e-29
+ drout = 8.376749865e-01 ldrout = 8.291329327e-8
+ pscbe1 = 1.037253098e+09 lpscbe1 = -3.066279457e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.174946640e-06 lalpha0 = -1.672796894e-12
+ alpha1 = 0.85
+ beta0 = 1.689804911e+01 lbeta0 = 5.720552343e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.702718609e-01 lkt1 = -4.432457430e-9
+ kt2 = -1.732617328e-02 lkt2 = -9.905380073e-9
+ at = 1.158432509e+05 lat = -5.372855313e-2
+ ute = -8.338566440e-01 lute = -2.433498184e-7
+ ua1 = 1.741162744e-09 lua1 = -4.645563804e-16
+ ub1 = -7.096737806e-19 lub1 = 3.973648481e-26
+ uc1 = 7.705161066e-11 luc1 = -3.642475369e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.150 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.316084900e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.980291269e-8
+ k1 = 2.425254334e-02 lk1 = 2.302273434e-7
+ k2 = 1.364915753e-01 lk2 = -7.397047947e-08 wk2 = -8.326672685e-23 pk2 = -2.081668171e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.555850181e-01 ldsub = 7.902988866e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
+ voff = {-1.072895691e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.856546771e-8
+ nfactor = 4.181852129e+00 lnfactor = -7.003856918e-7
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.461928472e-02 letab = -2.311014721e-08 wetab = 8.673617380e-24 petab = 2.168404345e-30
+ u0 = 1.451973038e-02 lu0 = 1.503840623e-9
+ ua = -2.102031242e-09 lua = 2.598939142e-16 wua = -3.308722450e-30
+ ub = 2.286030502e-18 lub = -3.339470352e-25
+ uc = 1.078724767e-11 luc = 2.132518899e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.752347497e+05 lvsat = -6.761528150e-4
+ a0 = 1.264221183e+00 la0 = 6.148781451e-8
+ ags = -9.846887499e-01 lags = 5.827755403e-07 wags = -4.440892099e-22 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.220181432e-02 lketa = -4.051305667e-08 wketa = 2.775557562e-23 pketa = 2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.742500265e-01 lpclm = -1.136192514e-7
+ pdiblc1 = -3.048846468e-01 lpdiblc1 = 1.726029866e-07 wpdiblc1 = -2.220446049e-22 ppdiblc1 = 5.551115123e-29
+ pdiblc2 = -8.673906560e-03 lpdiblc2 = 4.454229746e-09 wpdiblc2 = 3.361026735e-24 ppdiblc2 = -1.978668965e-30
+ pdiblcb = -8.553970447e-02 lpdiblcb = -4.630533306e-9
+ drout = 1.518101611e+00 ldrout = -2.646391004e-7
+ pscbe1 = 6.718076254e+07 lpscbe1 = 1.888714225e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.945729689e-06 lalpha0 = -2.066502085e-12
+ alpha1 = 0.85
+ beta0 = 2.187554651e+01 lbeta0 = -1.970380753e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.185774105e-01 lkt1 = 2.024134103e-8
+ kt2 = -4.489649533e-02 lkt2 = 4.177154445e-9
+ at = -8.189373154e+03 lat = 9.625574790e-3
+ ute = -1.301136473e+00 lute = -4.669823687e-9
+ ua1 = 1.724096898e-09 lua1 = -4.558393851e-16
+ ub1 = -2.029308260e-18 lub1 = 7.137873019e-25 wub1 = 1.540743956e-39
+ uc1 = -1.418079323e-10 luc1 = 7.536563684e-17 wuc1 = -9.047287950e-32 puc1 = 1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.151 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.910376278e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.685600016e-8
+ k1 = 9.070734895e-01 lk1 = 9.610978680e-17
+ k2 = -1.545831667e-01 lk2 = 1.937738201e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.456701426e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999995e-03 lcdscd = 1.016985107e-18
+ cit = 0.0
+ voff = {-9.930380979e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804193e-8
+ nfactor = 3.328469708e-01 lnfactor = 3.033809674e-7
+ eta0 = 2.586027983e-03 leta0 = -4.933778854e-10
+ etab = -4.399800002e-02 letab = 4.149791621e-18
+ u0 = 4.971157021e-03 lu0 = 3.993974876e-9
+ ua = -1.140127232e-09 lua = 9.042815314e-18
+ ub = -1.341759587e-19 lub = 2.972089268e-25
+ uc = 1.349581004e-10 luc = -1.105683100e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.255953955e+05 lvsat = 1.226909581e-2
+ a0 = 1.499999998e+00 la0 = 2.935962584e-16
+ ags = 1.250000000e+00 lags = 6.285816312e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.230652295e-08 lb0 = -1.103294889e-14
+ b1 = -2.897739533e-08 lb1 = 7.556899020e-15
+ keta = -2.361801760e-01 lketa = 3.990864906e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.002113030e-01 lpclm = -4.215378882e-8
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026290495e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347644218e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990363595e-18
+ drout = 5.033266586e-01 ldrout = 2.662119414e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629852295e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.294319198e-09 lalpha0 = 5.970517983e-15
+ alpha1 = 0.85
+ beta0 = 1.556519520e+01 lbeta0 = -3.247294746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.664260576e-01 lkt1 = 6.640998307e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.595168442e-18
+ at = -3.941737010e+04 lat = 1.776939920e-2
+ ute = -1.327992328e+00 lute = 2.333807174e-9
+ ua1 = -2.384733758e-11 lua1 = 3.009865197e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190619704e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.152 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.663494217e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.487564257e-09 wvth0 = 2.944699932e-08 pvth0 = -5.618075213e-15
+ k1 = 0.90707349
+ k2 = -1.642822690e-02 lk2 = -2.442029014e-08 wk2 = -2.380983222e-08 pk2 = 4.542582650e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.666911915e+00 ldsub = -4.213092735e-07 wdsub = -9.761079297e-07 pdsub = 1.862277275e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -2.079586503e-19
+ cit = 0.0
+ voff = {-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.724309667e-17
+ nfactor = -3.997892211e+00 lnfactor = 1.129625373e-06 wnfactor = 1.621326138e-06 pnfactor = -3.093263285e-13
+ eta0 = -1.264693740e-02 leta0 = 2.412858647e-09 weta0 = 3.944984598e-09 peta0 = -7.526478316e-16
+ etab = -0.043998
+ u0 = -1.293558438e-01 lu0 = 2.962168606e-08 wu0 = 5.846163092e-08 pu0 = -1.115366072e-14
+ ua = -1.023245120e-09 lua = -1.325665546e-17 wua = 1.329012897e-16 pua = -2.535570545e-23
+ ub = -4.555562994e-18 lub = 1.140747674e-24 wub = 5.016704073e-25 pub = -9.571169033e-32
+ uc = -2.367505281e-10 luc = 5.985997139e-17 wuc = 1.138127893e-16 puc = -2.171388681e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.842833836e+06 lvsat = -2.962773573e-01 wvsat = -6.372424012e-01 pvsat = 1.215769288e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.404690650e-06 lb0 = -6.525287670e-13 wb0 = -3.644673002e-13 pb0 = 6.953525834e-20
+ b1 = 2.645164180e-06 lb1 = -5.026318756e-13 wb1 = -1.372712398e-12 pb1 = 2.618943076e-19
+ keta = -8.680495464e-01 lketa = 1.604604788e-07 wketa = 3.716866934e-07 pketa = -7.091261748e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.238616222e-02 lpclm = 3.183781848e-08 wpclm = 1.113923637e-07 ppclm = -2.125210350e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000016e-08 lalpha0 = -2.923100113e-23 walpha0 = 2.103028225e-22 palpha0 = -4.012283898e-29
+ alpha1 = 0.85
+ beta0 = 1.393352521e+01 lbeta0 = -1.342968489e-08 wbeta0 = 3.808509064e-17 pbeta0 = -7.275957614e-24
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.815416658e-01 lkt1 = -9.553755267e-09 wkt1 = -7.824496606e-17 pkt1 = 1.492805879e-23
+ kt2 = -0.028878939
+ at = 5.372048689e+04 lat = 1.763598993e-11 wat = -2.483697608e-11 pat = 4.738511052e-18
+ ute = -1.159677081e+00 lute = -2.977838545e-08 wute = -2.128336404e-07 pute = 4.060567893e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.153 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.154 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.305913336e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.011998805e-06 wvth0 = 1.002040773e-08 pvth0 = -2.005162347e-13
+ k1 = 7.868894831e-01 lk1 = -4.379996120e-06 wk1 = -7.182648365e-08 pk1 = 1.437304393e-12
+ k2 = -1.195722482e-01 lk2 = 1.753665286e-06 wk2 = 3.054281727e-08 pk2 = -6.111857802e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.014231969e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.371667962e-07 wvoff = -9.655247898e-11 pvoff = 1.932090995e-15
+ nfactor = 4.776205409e+00 lnfactor = -1.708931949e-05 wnfactor = -1.724151410e-07 pnfactor = 3.450162491e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.586123952e-02 lu0 = 1.229274687e-07 wu0 = 1.508846931e-09 pu0 = -3.019321304e-14
+ ua = -1.567945616e-09 lua = 1.038160210e-14 wua = 1.362153298e-16 pua = -2.725775815e-21
+ ub = 1.305420030e-18 lub = -1.142016165e-24 wub = -5.318277982e-27 pub = 1.064229226e-31
+ uc = 6.333423789e-11 luc = -2.961043608e-16 wuc = 1.458237511e-20 puc = -2.918047878e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.116168035e+00 la0 = 4.931297306e-06 wa0 = 1.132278538e-07 pa0 = -2.265778352e-12
+ ags = 3.189492136e-01 lags = 5.188954170e-07 wags = 7.462744911e-10 pags = -1.493353914e-14
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.577685926e-08 lb0 = -8.020494973e-13 wb0 = -1.548761980e-14 pb0 = 3.099194454e-19
+ b1 = 1.533352558e-08 lb1 = -5.920242223e-14 wb1 = 7.533083426e-16 pb1 = -1.507429204e-20
+ keta = -4.819492937e-03 lketa = 5.460802153e-09 wketa = 8.927844716e-10 pketa = -1.786531901e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.567951267e-02 lpclm = -5.764009390e-07 wpclm = -2.286516418e-08 ppclm = 4.575499072e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 2.763457643e-03 lpdiblc2 = -3.608205223e-08 wpdiblc2 = -9.118428639e-10 ppdiblc2 = 1.824669241e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -1.004485635e+08 lpscbe1 = 6.512481558e+03 wpscbe1 = 1.031667870e+01 ppscbe1 = -2.064448497e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.979454292e-01 lkt1 = 2.314333279e-07 wkt1 = 6.073130341e-09 pkt1 = -1.215281116e-13
+ kt2 = -5.740837429e-02 lkt2 = 5.581096922e-07 wkt2 = 9.028723014e-09 pkt2 = -1.806718441e-13
+ at = 2.296000487e+05 lat = -1.092589891e+00 wat = -1.286680157e-02 pat = 2.574748127e-7
+ ute = -6.770835021e-01 lute = -8.771057639e-06 wute = -1.393903503e-07 pute = 2.789310471e-12
+ ua1 = 1.509250306e-09 lua1 = -7.769193781e-15 wua1 = -1.976340721e-16 pua1 = 3.954813123e-21
+ ub1 = -8.022631173e-19 lub1 = 4.658373252e-24 wub1 = 1.731785713e-25 pub1 = -3.465439329e-30
+ uc1 = 1.513892071e-10 luc1 = -2.352685020e-15 wuc1 = -3.374747090e-17 puc1 = 6.753134183e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.155 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.251093781e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.548349776e-07 wvth0 = -9.063576713e-09 pvth0 = -4.763851928e-14
+ k1 = -9.731408218e-02 lk1 = 2.703169421e-06 wk1 = 2.198486255e-07 pk1 = -8.992424877e-13
+ k2 = 2.511914443e-01 lk2 = -1.216443311e-06 wk2 = -9.485651157e-08 pk2 = 3.933614077e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.283237652e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.059860198e-07 wvoff = -1.036592696e-08 pvoff = 8.419785228e-14
+ nfactor = 3.799359222e+00 lnfactor = -9.264013724e-06 wnfactor = 8.042150399e-08 pnfactor = 1.424742234e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.111833772e-02 lu0 = 7.061200158e-10 wu0 = -3.050535332e-09 pu0 = 6.331022559e-15
+ ua = -1.238479865e-10 lua = -1.186754974e-15 wua = -3.504206920e-16 pua = 1.172561216e-21
+ ub = 9.800139738e-19 lub = 1.464742117e-24 wub = 1.532480793e-25 pub = -1.163818232e-30
+ uc = -6.280647041e-11 luc = 7.143818593e-16 wuc = 2.976625492e-17 puc = -2.386260867e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.047189575e+00 la0 = -2.526917007e-06 wa0 = -2.623788062e-07 pa0 = 7.431262215e-13
+ ags = 2.172567339e-01 lags = 1.333532110e-06 wags = 5.912826808e-08 pags = -4.826191961e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.729213055e-07 lb0 = 7.896789789e-13 wb0 = 7.069918857e-14 pb0 = -3.805046325e-19
+ b1 = 1.474336057e-08 lb1 = -5.447473666e-14 wb1 = -3.564313932e-15 pb1 = 1.951325603e-20
+ keta = -1.198656708e-02 lketa = 6.287469937e-08 wketa = -2.292473845e-09 pketa = 7.651103722e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.799318387e+00 lpclm = 1.420348241e-05 wpclm = 4.523878342e-07 ppclm = -3.349600158e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -3.516886206e-03 lpdiblc2 = 1.422843835e-08 wpdiblc2 = 7.602127475e-10 ppdiblc2 = 4.852212732e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 9.915650021e+08 lpscbe1 = -2.235405425e+03 wpscbe1 = -1.453572731e+02 ppscbe1 = 1.040625864e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.975461713e-01 lkt1 = 2.282349584e-07 wkt1 = 4.662816536e-09 pkt1 = -1.102303895e-13
+ kt2 = 1.762431711e-02 lkt2 = -4.296114161e-08 wkt2 = -1.125627331e-08 pkt2 = -1.817307950e-14
+ at = 4.629423130e+04 lat = 3.758337852e-01 wat = 3.860040471e-02 pat = -1.548179628e-7
+ ute = -2.561128647e+00 lute = 6.321624833e-06 wute = 5.480430399e-07 pute = -2.717571307e-12
+ ua1 = -1.235537772e-09 lua1 = 1.421871612e-14 wua1 = 1.134331838e-15 pua1 = -6.715280743e-21
+ ub1 = 1.045270910e-18 lub1 = -1.014182647e-23 wub1 = -8.544585660e-25 pub1 = 4.766741863e-30
+ uc1 = -2.568724225e-10 luc1 = 9.178115262e-16 wuc1 = 7.629790755e-17 puc1 = -2.062365587e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.156 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.449600164e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.258602848e-07 wvth0 = -4.210660109e-08 pvth0 = 8.488998031e-14
+ k1 = 6.767922676e-01 lk1 = -4.016054889e-07 wk1 = -4.851042420e-08 pk1 = 1.770882319e-13
+ k2 = -1.140809945e-01 lk2 = 2.485862726e-07 wk2 = 2.836213145e-08 pk2 = -1.008422007e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.802460648e+00 ldsub = -4.983243772e-06 wdsub = -3.875632348e-07 pdsub = 1.554433196e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.185389296e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.981960633e-07 wvoff = 3.335381783e-08 pvoff = -9.115268803e-14
+ nfactor = -1.302471700e+00 lnfactor = 1.119833831e-05 wnfactor = 1.308493788e-06 pnfactor = -3.500792888e-12
+ eta0 = 4.092520717e-01 leta0 = -1.320559600e-06 weta0 = -1.027042572e-07 peta0 = 4.119247970e-13
+ etab = -3.578367167e-01 letab = 1.154451474e-06 wetab = 8.978548273e-08 petab = -3.601103571e-13
+ u0 = 3.292302386e-02 lu0 = -6.532089871e-09 wu0 = -1.390777024e-09 pu0 = -3.259128268e-16
+ ua = -1.372457982e-09 lua = 3.821152515e-15 wua = 2.743738166e-16 pua = -1.333355852e-21
+ ub = 3.374251416e-18 lub = -8.138031897e-24 wub = -7.791033910e-25 pub = 2.575643992e-30
+ uc = 1.634440429e-10 luc = -1.930605318e-16 wuc = -5.272783789e-17 puc = 9.224006587e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.932576895e+05 lvsat = -8.553309555e-01 wvsat = -8.784766655e-02 pvsat = 3.523381911e-7
+ a0 = 4.047405694e+00 la0 = -1.054935582e-05 wa0 = -1.001047615e-06 pa0 = 3.705768740e-12
+ ags = -2.910547498e-02 lags = 2.321638208e-06 wags = 1.460667578e-07 pags = -8.313108734e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.094130473e-07 lb0 = 9.360395460e-13 wb0 = 6.545155449e-14 pb0 = -3.594574952e-19
+ b1 = -1.774042840e-08 lb1 = 7.581078938e-14 wb1 = 4.510421413e-15 pb1 = -1.287277944e-20
+ keta = 4.282352676e-02 lketa = -1.569568577e-07 wketa = -1.744319475e-08 pketa = 6.841740302e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.036177216e+00 lpclm = -2.123379966e-05 wpclm = -2.436380297e-06 ppclm = 8.236630620e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.239717606e-02 lpdiblc2 = -4.959945979e-08 wpdiblc2 = -4.104489560e-09 ppdiblc2 = 2.436349264e-14
+ pdiblcb = -7.676919366e-02 lpdiblcb = 2.076351572e-07 wpdiblcb = 1.614846812e-08 ppdiblcb = -6.476804984e-14
+ drout = 0.56
+ pscbe1 = 6.646040177e+07 lpscbe1 = 1.474991155e+03 wpscbe1 = 2.288144740e+02 ppscbe1 = -4.600969408e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.099213957e-01 lkt1 = -5.242878645e-07 wkt1 = -6.102148779e-08 pkt1 = 1.532152987e-13
+ kt2 = 1.182831932e-01 lkt2 = -4.466823525e-07 wkt2 = -5.468480051e-08 pkt2 = 1.560094494e-13
+ at = 2.668552321e+05 lat = -5.087891891e-01 wat = -3.957020627e-02 pat = 1.587076293e-7
+ ute = 1.475554346e+00 lute = -9.868646804e-06 wute = -9.645923141e-07 pute = 3.349285394e-12
+ ua1 = 9.963154521e-09 lua1 = -3.069684215e-14 wua1 = -3.214224497e-15 pua1 = 1.072584813e-20
+ ub1 = -6.397255323e-18 lub1 = 1.970855355e-23 wub1 = 2.017183453e-24 pub1 = -6.750799742e-30
+ uc1 = -1.487316875e-10 luc1 = 4.840821802e-16 wuc1 = 6.456176813e-17 puc1 = -1.591654151e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.157 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.416120062e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.830290472e-07 wvth0 = 2.039514383e-08 pvth0 = -4.078765335e-14
+ k1 = 4.982244104e-01 lk1 = -4.254374149e-08 wk1 = 3.871683499e-08 pk1 = 1.692880326e-15
+ k2 = 2.288641947e-02 lk2 = -2.682588582e-08 wk2 = -2.723736238e-08 pk2 = 1.095648308e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.621685496e+00 ldsub = 1.901981355e-06 wdsub = 7.751264696e-07 pdsub = -7.834869837e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {4.248839559e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.266740278e-07 wvoff = -4.369677986e-08 pvoff = 6.377957509e-14
+ nfactor = 7.381643048e+00 lnfactor = -6.263558046e-06 wnfactor = -1.300748206e-06 pnfactor = 1.745834383e-12
+ eta0 = -5.001998154e-01 leta0 = 5.081535227e-07 weta0 = 2.054085144e-07 peta0 = -2.076240507e-13
+ etab = 7.852496013e-01 letab = -1.144050491e-06 wetab = -2.887519434e-07 petab = 4.010473998e-13
+ u0 = 3.018844128e-02 lu0 = -1.033429503e-09 wu0 = -1.417053343e-10 pu0 = -2.837528693e-15
+ ua = 1.933638684e-09 lua = -2.826700375e-15 wua = -6.730837394e-16 pua = 5.717785370e-22
+ ub = -2.915551493e-18 lub = 4.509415736e-24 wub = 1.080273374e-24 pub = -1.163164776e-30
+ uc = 1.050319021e-10 luc = -7.560621687e-17 wuc = -1.766516822e-17 puc = 2.173654055e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -5.805411377e+04 lvsat = -1.489180998e-01 wvsat = 5.544656986e-02 pvsat = 6.420414669e-8
+ a0 = -2.677942814e+00 la0 = 2.973880810e-06 wa0 = 1.303234058e-06 pa0 = -9.276485887e-13
+ ags = -2.303825178e+00 lags = 6.895612740e-06 wags = 8.231973570e-07 pags = -2.192875602e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.447998951e-07 lb0 = 1.811509324e-12 wb0 = 2.423431492e-13 pb0 = -7.151486374e-19
+ b1 = -1.808193556e-08 lb1 = 7.649748719e-14 wb1 = 7.400223458e-15 pb1 = -1.868355294e-20
+ keta = 2.462311287e-01 lketa = -5.659660159e-07 wketa = -7.117456941e-08 pketa = 1.764596990e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.444852107e+00 lpclm = 7.884451368e-06 wpclm = 3.123210116e-06 ppclm = -2.942515948e-12
+ pdiblc1 = 1.167079867e+00 lpdiblc1 = -1.562541318e-06 wpdiblc1 = -3.052679362e-07 ppdiblc1 = 6.138284924e-13
+ pdiblc2 = -2.581068363e-02 lpdiblc2 = 2.722836956e-08 wpdiblc2 = 1.462482297e-08 ppdiblc2 = -1.329714678e-14
+ pdiblcb = -2.475802147e-02 lpdiblcb = 1.030518203e-07 wpdiblcb = -7.548084717e-11 ppdiblcb = -3.214516040e-14
+ drout = -6.406317959e-01 ldrout = 2.414213606e-06 wdrout = 3.448070684e-07 pdrout = -6.933332258e-13
+ pscbe1 = 1.075235807e+09 lpscbe1 = -5.534403071e+02 wpscbe1 = -8.585485570e+01 ppscbe1 = 1.726357419e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.282899291e-05 lalpha0 = 4.596454292e-11 walpha0 = 7.130451377e-12 palpha0 = -1.433781180e-17
+ alpha1 = 0.85
+ beta0 = -1.146158552e+00 lbeta0 = 3.017417353e-05 wbeta0 = 4.680901049e-06 pbeta0 = -9.412290297e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.349159301e-01 lkt1 = 3.302851953e-07 wkt1 = 5.820385706e-08 pkt1 = -8.652135556e-14
+ kt2 = -1.793184377e-01 lkt2 = 1.517308404e-07 wkt2 = 4.518360462e-08 pkt2 = -4.480454149e-14
+ at = 1.766676771e+05 lat = -3.274413161e-01 wat = -8.284856880e-03 pat = 9.579948677e-8
+ ute = -4.694601147e+00 lute = 2.538215479e-06 wute = 9.479945560e-07 pute = -4.965175086e-13
+ ua1 = -9.080467514e-09 lua1 = 7.595806433e-15 wua1 = 3.077194516e-15 pua1 = -1.924849145e-21
+ ub1 = 5.339270394e-18 lub1 = -3.891088049e-24 wub1 = -1.795278181e-24 pub1 = 9.152447362e-31
+ uc1 = 1.641971944e-10 luc1 = -1.451508344e-16 wuc1 = -3.784801648e-17 puc1 = 4.675874607e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.158 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.049961088e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.788268370e-08 wvth0 = -2.049622307e-08 pvth0 = 5.447678252e-16
+ k1 = 7.571772566e-01 lk1 = -3.042896532e-07 wk1 = -5.028662417e-08 pk1 = 9.165633079e-14
+ k2 = -1.151727407e-01 lk2 = 1.127223804e-07 wk2 = 1.475527961e-08 pk2 = -3.148909155e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.924073019e-01 ldsub = 6.832175295e-08 wdsub = 6.673439569e-09 pdsub = -6.745419288e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-3.146488068e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.343152565e-07 wvoff = 7.791534794e-08 pvoff = -5.914426111e-14
+ nfactor = -4.064411422e+00 lnfactor = 5.305953568e-06 wnfactor = 2.340341541e-06 pnfactor = -1.934528158e-12
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 2.688821388e-23 peta0 = 2.818925648e-29
+ etab = -6.990280776e-01 letab = 3.562366066e-07 wetab = 2.179517475e-07 petab = -1.111215972e-13
+ u0 = 4.827238984e-02 lu0 = -1.931243154e-08 wu0 = -8.907568867e-09 pu0 = 6.022883444e-15
+ ua = 1.278271205e-09 lua = -2.164264102e-15 wua = -7.918139063e-16 pua = 6.917893275e-22
+ ub = -2.326669368e-19 lub = 1.797593587e-24 wub = 5.537067210e-25 pub = -6.309185751e-31
+ uc = -1.459348637e-10 luc = 1.780674764e-16 wuc = 7.094448321e-17 puc = -6.782885457e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.403778985e+05 lvsat = 7.429224293e-01 wvsat = 3.415697057e-01 pvsat = -2.250051133e-7
+ a0 = -5.126263919e-01 la0 = 7.852092845e-07 wa0 = 6.278025757e-07 pa0 = -2.449319025e-13
+ ags = 8.538587052e+00 lags = -4.063745747e-06 wags = -2.542132338e-06 pags = 1.208752539e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.860318738e-06 lb0 = -7.206295186e-13 wb0 = -7.512278901e-13 pb0 = 2.891390592e-19
+ b1 = 1.576279736e-07 lb1 = -1.011076291e-13 wb1 = -3.937323738e-14 pb1 = 2.859440645e-20
+ keta = -6.098014576e-01 lketa = 2.992997378e-07 wketa = 2.019950221e-07 pketa = -9.965629978e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.967141068e-01 lpclm = -4.460083784e-07 wpclm = 2.064539015e-07 ppclm = 5.700398618e-15
+ pdiblc1 = 6.875439659e-01 lpdiblc1 = -1.077833142e-06 wpdiblc1 = -2.021418899e-09 ppdiblc1 = 3.073111581e-13
+ pdiblc2 = 6.305515001e-03 lpdiblc2 = -5.234234385e-09 wpdiblc2 = 1.292475416e-09 ppdiblc2 = 1.790034709e-16
+ pdiblcb = 4.745042074e-01 lpdiblcb = -4.015954510e-07 wpdiblcb = -1.558113464e-07 ppdiblcb = 1.252704722e-13
+ drout = 2.511772333e+00 ldrout = -7.721923531e-07 wdrout = -6.896142680e-07 pdrout = 3.522453791e-13
+ pscbe1 = 1.777321433e+09 lpscbe1 = -1.263098629e+03 wpscbe1 = -3.048578294e+02 ppscbe1 = 3.940008816e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.127868928e-05 lalpha0 = -8.726744729e-12 walpha0 = -9.929102912e-12 palpha0 = 2.905746839e-18
+ alpha1 = 0.85
+ beta0 = 3.191939782e+01 lbeta0 = -3.248027931e-06 wbeta0 = -6.187774215e-06 pbeta0 = 1.573614498e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.214628087e-01 lkt1 = 1.345116850e-08 wkt1 = -2.010601048e-08 pkt1 = -7.366837796e-15
+ kt2 = -6.347895933e-02 lkt2 = 3.464191743e-08 wkt2 = 1.901180946e-08 pkt2 = -1.835045736e-14
+ at = -3.425754759e+05 lat = 1.974023935e-01 wat = 1.888373430e-01 pat = -1.034488731e-7
+ ute = -3.630682652e+00 lute = 1.462821559e-06 wute = 1.152102131e-06 pute = -7.028265880e-13
+ ua1 = -5.458360167e-09 lua1 = 3.934631036e-15 wua1 = 2.965713872e-15 pua1 = -1.812166071e-21
+ ub1 = 5.839485692e-18 lub1 = -4.396698668e-24 wub1 = -2.697808360e-24 pub1 = 1.827509606e-30
+ uc1 = 3.562791845e-10 luc1 = -3.393046209e-16 wuc1 = -1.150227729e-16 puc1 = 1.247659095e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.159 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {7.279779487e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.493471836e-08 wvth0 = -3.969766388e-08 pvth0 = 1.035259497e-14
+ k1 = -6.163447123e-01 lk1 = 3.972861393e-07 wk1 = 2.638825087e-07 pk1 = -6.881686392e-14
+ k2 = 3.690765777e-01 lk2 = -1.346253919e-07 wk2 = -9.580920520e-08 pk2 = 2.498569939e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.879857035e-01 ldsub = 7.058024352e-08 wdsub = -1.334687914e-08 pdsub = 3.480679223e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446113e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
+ voff = {8.056854541e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.755623395e-08 wvoff = -7.738476881e-08 pvoff = 2.018086432e-14
+ nfactor = 1.135890527e+01 lnfactor = -2.572060672e-06 wnfactor = -2.956457855e-06 pnfactor = 7.710028181e-13
+ eta0 = 1.000416472e+00 leta0 = -2.607135881e-7
+ etab = 4.262765349e-02 letab = -2.259075767e-08 wetab = 8.204166366e-10 petab = -2.139531730e-16
+ u0 = 2.161853998e-04 lu0 = 5.234004905e-09 wu0 = 5.892087891e-09 pu0 = -1.536574033e-15
+ ua = -4.892218647e-09 lua = 9.875357269e-16 wua = 1.149367478e-15 pua = -2.997389472e-22
+ ub = 5.666131430e-18 lub = -1.215430036e-24 wub = -1.392371736e-24 pub = 3.631110555e-31
+ uc = 3.175505559e-10 luc = -5.867438711e-17 wuc = -1.263656231e-16 puc = 3.295438538e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.659573895e+05 lvsat = -1.286497472e-01 wvsat = -2.021443585e-01 pvsat = 5.271641867e-8
+ a0 = 5.287516015e-01 la0 = 2.532879847e-07 wa0 = 3.029634556e-07 pa0 = -7.900862772e-14
+ ags = -1.133500860e-01 lags = 3.555426155e-07 wags = -3.589322785e-07 pags = 9.360451319e-14
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.183809937e-07 lb0 = -2.395009058e-13 wb0 = -3.783105195e-13 pb0 = 9.865808713e-20
+ b1 = -8.237386775e-08 lb1 = 2.148195148e-14 wb1 = 3.393243209e-14 pb1 = -8.849103235e-21
+ keta = 3.802209938e-02 lketa = -3.159946554e-08 wketa = 1.407971833e-08 pketa = -3.671793425e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -4.050947308e-01 lpclm = 1.678587505e-07 wpclm = 4.446166446e-07 ppclm = -1.159497963e-13
+ pdiblc1 = -3.278954597e+00 lpdiblc1 = 9.481987926e-07 wpdiblc1 = 1.225114583e-06 ppdiblc1 = -3.194927315e-13
+ pdiblc2 = -1.682264780e-02 lpdiblc2 = 6.579307378e-09 wpdiblc2 = 3.356727276e-09 ppdiblc2 = -8.753874793e-16
+ pdiblcb = -5.291490169e-01 lpdiblcb = 1.110565648e-07 wpdiblcb = 1.827368713e-07 ppdiblcb = -4.765521772e-14
+ drout = 1.518100973e+00 ldrout = -2.646389342e-07 wdrout = 2.625333235e-13 pdrout = -6.846501532e-20
+ pscbe1 = -2.246635793e+09 lpscbe1 = 7.922823868e+02 wpscbe1 = 9.531350815e+02 ppscbe1 = -2.485642854e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.897735550e-05 lalpha0 = -7.551255653e-12 walpha0 = -8.663599683e-12 palpha0 = 2.259345507e-18
+ alpha1 = 0.85
+ beta0 = 3.728599233e+01 lbeta0 = -5.989209276e-06 wbeta0 = -6.348055768e-06 pbeta0 = 1.655484071e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.473189847e-01 lkt1 = -2.442045880e-08 wkt1 = -7.054682586e-08 pkt1 = 1.839762453e-14
+ kt2 = 3.899590679e-02 lkt2 = -1.770080953e-08 wkt2 = -3.455796499e-08 pkt2 = 9.012233458e-15
+ at = 5.971894237e+04 lat = -8.083963181e-03 wat = -2.797360823e-02 pat = 7.295125396e-9
+ ute = -1.907692392e-01 lute = -2.942380531e-07 wute = -4.573957954e-07 pute = 1.192824199e-13
+ ua1 = 4.611184524e-09 lua1 = -1.208751419e-15 wua1 = -1.189283780e-15 pua1 = 3.101485598e-22
+ ub1 = -6.394172991e-18 lub1 = 1.852082916e-24 wub1 = 1.798027458e-24 pub1 = -4.689003888e-31
+ uc1 = -7.828252591e-10 luc1 = 2.425339814e-16 wuc1 = 2.640555494e-16 puc1 = -6.886199051e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.160 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {-3.179394558e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.532031549e-07 wvth0 = 2.153710557e-07 pvth0 = -5.616575613e-14
+ k1 = 9.070734895e-01 lk1 = 9.610845453e-17
+ k2 = -2.578321670e-01 lk2 = 2.886363201e-08 wk2 = 4.253156721e-08 pk2 = -1.109163729e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.862269127e+00 ldsub = -3.660494333e-07 wdsub = -5.782038727e-07 pdsub = 1.507874752e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999993e-03 lcdscd = 1.467913464e-18 wcdscd = 7.122653162e-19 pcdscd = -1.857489856e-25
+ cit = 0.0
+ voff = {-9.930380956e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.064804199e-08 wvoff = -9.330769490e-17 pvoff = 2.433334090e-23
+ nfactor = -1.228664795e+01 lnfactor = 3.594368570e-06 wnfactor = 5.198373782e-06 pnfactor = -1.355663105e-12
+ eta0 = 2.586026044e-03 leta0 = -4.933773123e-10 weta0 = 9.052863693e-16 peta0 = -2.360860111e-22
+ etab = -4.399800002e-02 letab = 4.149736110e-18
+ u0 = -3.673397487e-02 lu0 = 1.487008940e-08 wu0 = 1.717967839e-08 pu0 = -4.480219608e-15
+ ua = -1.206504277e-09 lua = 2.635301933e-17 wua = 2.734282884e-17 pua = -7.130626962e-24
+ ub = -2.283224180e-18 lub = 8.576506162e-25 wub = 8.852617319e-25 pub = -2.308638660e-31
+ uc = 2.578509145e-10 luc = -4.310555642e-17 wuc = -5.062348271e-17 puc = 1.320189556e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.212823632e+04 lvsat = 9.512697086e-02 wvsat = 1.308805311e-01 pvsat = -3.413181018e-8
+ a0 = 1.499999998e+00 la0 = 2.935935939e-16
+ ags = 1.250000000e+00 lags = 6.286082765e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.239601204e-07 lb0 = 1.105628639e-13 wb0 = 1.920701509e-13 pb0 = -5.008920638e-20
+ b1 = -4.775969536e-07 lb1 = 1.245505991e-13 wb1 = 1.848007519e-13 pb1 = -4.819344888e-20
+ keta = -5.879486345e-01 lketa = 1.316449383e-07 wketa = 1.449046846e-07 pketa = -3.778911308e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.162516963e-01 lpclm = -4.633689883e-08 wpclm = -6.607551306e-09 ppclm = 1.723156875e-15
+ pdiblc1 = 3.569721503e-01 lpdiblc1 = -5.026246086e-17
+ pdiblc2 = 8.406112093e-03 lpdiblc2 = 1.347651157e-18
+ pdiblcb = -1.032957700e-01 lpdiblcb = 3.990363595e-18
+ drout = 5.033266586e-01 ldrout = 2.662110532e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 2.629947662e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.823435072e-07 lalpha0 = -4.191965620e-14 walpha0 = -7.564629709e-14 palpha0 = 1.972749523e-20
+ alpha1 = 0.85
+ beta0 = 2.012949758e+01 lbeta0 = -1.515035635e-06 wbeta0 = -1.880182208e-06 pbeta0 = 4.903251974e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.758255074e-01 lkt1 = -1.698635676e-08 wkt1 = -3.732126582e-08 pkt1 = 9.732863628e-15
+ kt2 = -2.887893901e-02 lkt2 = 1.595196197e-18
+ at = -1.244348822e+05 lat = 3.994077611e-02 wat = 3.502143379e-02 pat = -9.133099632e-9
+ ute = -1.015837471e+00 lute = -7.907180915e-08 wute = -1.285865742e-07 pute = 3.353357834e-14
+ ua1 = -2.384733758e-11 lua1 = 3.009865455e-25
+ ub1 = 7.077531678e-19 lub1 = 4.275656921e-34
+ uc1 = 1.471862500e-10 luc1 = -6.190878198e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.161 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {1.239660536e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.937255989e-08 wvth0 = -2.479113947e-07 pvth0 = 3.222204945e-14
+ k1 = 0.90707349
+ k2 = 6.024711742e-02 lk2 = -3.182144236e-08 wk2 = -5.539486016e-08 pk2 = 7.591354085e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -7.208291699e-01 ldsub = 1.267695583e-07 wdsub = 4.194110310e-07 pdsub = -3.954348187e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000005e-03 lcdscd = -8.566584941e-19 wcdscd = -1.661955296e-18 pcdscd = 2.672189726e-25
+ cit = 0.0
+ voff = {-2.075300007e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.122231197e-16 wvoff = 2.177178438e-16 pvoff = -3.500599810e-23
+ nfactor = 2.544759612e+01 lnfactor = -3.604796918e-06 wnfactor = -1.050821276e-05 pnfactor = 1.640933715e-12
+ eta0 = -1.264693491e-02 leta0 = 2.412858568e-09 weta0 = 3.944984094e-09 peta0 = -7.526477988e-16
+ etab = -0.043998
+ u0 = 1.596124794e-01 lu0 = -2.259006522e-08 wu0 = -6.057366839e-08 pu0 = 1.035403041e-14
+ ua = -8.683663778e-10 lua = -3.815895797e-17 wua = 6.910177977e-17 pua = -1.509765017e-23
+ ub = 4.588753830e-19 lub = 3.344964090e-25 wub = -1.563937222e-24 pub = 2.364090056e-31
+ uc = -5.103733979e-10 luc = 1.034608872e-16 wuc = 2.265268053e-16 puc = -3.967449928e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.098033487e+05 lvsat = -3.879174852e-02 wvsat = -1.293176865e-01 pvsat = 1.551036697e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.492642732e-06 lb0 = -8.274561278e-13 wb0 = -8.126295770e-13 pb0 = 1.415934359e-19
+ b1 = 3.691851968e-06 lb1 = -6.709218828e-13 wb1 = -1.803876592e-12 pb1 = 3.312183469e-19
+ keta = -4.725592225e-02 lketa = 2.848833847e-08 wketa = 3.357553419e-08 pketa = -1.654906979e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.504117521e-02 lpclm = 3.785560295e-08 wpclm = 1.268098817e-07 ppclm = -2.373102149e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.984882588e-07 lalpha0 = 6.889491310e-14 walpha0 = 1.765080257e-13 palpha0 = -2.838001940e-20
+ alpha1 = 0.85
+ beta0 = 3.283486342e+00 lbeta0 = 1.698947464e-06 wbeta0 = 4.387091812e-06 pbeta0 = -7.053829438e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.929429503e-01 lkt1 = 2.443661169e-08 wkt1 = 8.708295386e-08 pkt1 = -1.400171983e-14
+ kt2 = -0.028878939
+ at = 2.520946815e+05 lat = -3.189579323e-02 wat = -8.171667875e-02 pat = 1.313889791e-8
+ ute = -1.912586392e+00 lute = 9.201533043e-08 wute = 9.731379786e-08 pute = -9.565050043e-15
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.162 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.163 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.627150263e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.691784641e-7
+ k1 = 5.566262089e-01 lk1 = 2.277529835e-7
+ k2 = -2.165726269e-02 lk2 = -2.056905354e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017327274e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.309728469e-7
+ nfactor = 4.223472310e+00 lnfactor = -6.028695726e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.069834161e-02 lu0 = 2.613325382e-8
+ ua = -1.131262846e-09 lua = 1.643236638e-15
+ ub = 1.288370552e-18 lub = -8.008426962e-25
+ uc = 6.338098646e-11 luc = -2.970398364e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.479156936e+00 la0 = -2.332395909e-6
+ ags = 3.213416405e-01 lags = 4.710210753e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.387376907e-08 lb0 = 1.914986009e-13
+ b1 = 1.774850174e-08 lb1 = -1.075279933e-13
+ keta = -1.957380452e-03 lketa = -5.181231829e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.762224597e-02 lpclm = 8.904248667e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.597527482e-04 lpdiblc2 = 2.241368535e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -6.737507727e+07 lpscbe1 = 5.850655103e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.784760245e-01 lkt1 = -1.581647627e-7
+ kt2 = -2.846385108e-02 lkt2 = -2.109296763e-8
+ at = 1.883513100e+05 lat = -2.671702072e-01 wat = 1.164153218e-16
+ ute = -1.123944838e+00 lute = 1.709889326e-7
+ ua1 = 8.756696787e-10 lua1 = 4.909252558e-15
+ ub1 = -2.470825931e-19 lub1 = -6.451225409e-24
+ uc1 = 4.320065665e-11 luc1 = -1.877470904e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.164 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.960531199e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.021141305e-7
+ k1 = 6.074825579e-01 lk1 = -1.796463452e-7
+ k2 = -5.290211314e-02 lk2 = 4.460527524e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.260637441e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.393772087e-8
+ nfactor = 4.057176644e+00 lnfactor = -4.696536728e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.133884946e-02 lu0 = 2.100228251e-8
+ ua = -1.247236071e-09 lua = 2.572273326e-15
+ ub = 1.471300791e-18 lub = -2.266257692e-24
+ uc = 3.261899065e-11 luc = -5.061207102e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.206048537e+00 la0 = -1.445829675e-7
+ ags = 4.068117269e-01 lags = -2.136614964e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.372805585e-08 lb0 = -4.301530117e-13 wb0 = 3.541366997e-30 pb0 = -3.319062208e-35
+ b1 = 3.316787051e-09 lb1 = 8.081384646e-15
+ keta = -1.933584143e-02 lketa = 8.740281358e-08 pketa = -2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.490412944e-01 lpclm = 3.465244080e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -1.079775722e-03 lpdiblc2 = 2.978379250e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.255747443e+08 lpscbe1 = 1.100660974e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.825979885e-01 lkt1 = -1.251445908e-7
+ kt2 = -1.846134680e-02 lkt2 = -1.012208889e-7
+ at = 1.700404475e+05 lat = -1.204858063e-1
+ ute = -8.041975216e-01 lute = -2.390438396e-6
+ ua1 = 2.400933761e-09 lua1 = -7.309311599e-15
+ ub1 = -1.693975356e-18 lub1 = 5.139522876e-24 pub1 = 3.081487911e-45
+ uc1 = -1.227453723e-11 luc1 = 2.566528161e-16 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.165 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.099735415e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.628229852e-8
+ k1 = 5.212762443e-01 lk1 = 1.661087306e-7
+ k2 = -2.315691021e-02 lk2 = -7.469636824e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.116123628e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.976323031e-9
+ nfactor = 2.892332897e+00 lnfactor = -2.459773863e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.846443345e-02 lu0 = -7.576909981e-9
+ ua = -4.928630170e-10 lua = -4.533555576e-16
+ ub = 8.765807986e-19 lub = 1.190369253e-25
+ uc = -5.592278815e-12 luc = 1.026451536e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.163327600e+04 lvsat = 2.742042995e-1
+ a0 = 8.382203100e-01 la0 = 1.330697336e-6
+ ags = 4.391592679e-01 lags = -3.434005609e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.133074850e-10 lb0 = -2.163189654e-13
+ b1 = -3.280798056e-09 lb1 = 3.454288663e-14
+ keta = -1.309633638e-02 lketa = 6.237749411e-08 wketa = 1.734723476e-24 pketa = -6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.744363068e-01 lpclm = 5.171412440e-06 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -7.611070267e-04 lpdiblc2 = 2.850568056e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.055457235e-01 lkt1 = -3.310613675e-8
+ kt2 = -5.702681193e-02 lkt2 = 5.345693870e-8
+ at = 140000.0
+ ute = -1.616761652e+00 lute = 8.685824428e-7
+ ua1 = -3.410928692e-10 lua1 = 3.688370421e-15
+ ub1 = 6.948567385e-20 lub1 = -1.933341932e-24
+ uc1 = 5.824216620e-11 luc1 = -2.617459078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.166 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.069953072e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.227089047e-8
+ k1 = 6.223438819e-01 lk1 = -3.711666019e-8
+ k2 = -6.443184982e-02 lk2 = 8.298702475e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.759591720e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.220774955e-8
+ nfactor = 3.211669446e+00 lnfactor = -6.667151992e-7
+ eta0 = 1.583043279e-01 leta0 = -1.574532464e-7
+ etab = -1.404391494e-01 letab = 1.416380554e-7
+ u0 = 2.973415850e-02 lu0 = -1.013005535e-8
+ ua = -2.241512811e-10 lua = -9.936773541e-16
+ ub = 5.476179603e-19 lub = 7.805107952e-25
+ uc = 4.840043040e-11 luc = -5.922630220e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.196979920e+05 lvsat = 5.690928146e-2
+ a0 = 1.5
+ ags = 3.352030625e-01 lags = -1.343668785e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.321102943e-07 lb0 = -4.811334227e-13 pb0 = -1.058791184e-34
+ b1 = 5.641899952e-09 lb1 = 1.660125039e-14
+ keta = 1.805777867e-02 lketa = -2.667642893e-10
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.567618932e+00 lpclm = -1.548745445e-6
+ pdiblc1 = 1.884437022e-01 lpdiblc1 = 4.052865819e-7
+ pdiblc2 = 2.107396742e-02 lpdiblc2 = -1.539998143e-8
+ pdiblcb = -0.025
+ drout = 4.647599830e-01 ldrout = 1.915072929e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.483244388e-01 lkt1 = 5.291270522e-8
+ kt2 = -3.446762206e-02 lkt2 = 8.095235534e-9
+ at = 1.501078600e+05 lat = -2.032474338e-2
+ ute = -1.655494688e+00 lute = 9.464662882e-7
+ ua1 = 7.844854756e-10 lua1 = 1.425073244e-15
+ ub1 = -4.160807111e-19 lub1 = -9.569718432e-25
+ uc1 = 4.286300461e-11 luc1 = 4.749612046e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.167 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.392887653e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.962911505e-8
+ k1 = 5.959670436e-01 lk1 = -1.045532135e-8
+ k2 = -6.786986822e-02 lk2 = 1.177380334e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.138011941e-01 ldsub = 4.669710627e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.486568763e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.529100738e-8
+ nfactor = 3.438318471e+00 lnfactor = -8.958088615e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = 1.214306433e-23 peta0 = 7.372574773e-29
+ etab = -0.0003125
+ u0 = 1.971626586e-02 lu0 = -4.109710889e-12
+ ua = -1.260147125e-09 lua = 5.349274039e-17
+ ub = 1.542420970e-18 lub = -2.250221600e-25
+ uc = 8.150086973e-11 luc = -3.938009089e-17 wuc = -5.169878828e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.546354561e+05 lvsat = 2.159498183e-2
+ a0 = 1.5
+ ags = 3.889507903e-01 lags = -1.886943293e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.479878483e-07 lb0 = 2.063002585e-13
+ b1 = 3.140418965e-08 lb1 = -9.438911366e-15
+ keta = 3.775962016e-02 lketa = -2.018110984e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.458569580e+00 lpclm = -4.277338871e-07 wpclm = -8.881784197e-22
+ pdiblc1 = 6.810636468e-01 lpdiblc1 = -9.264676145e-8
+ pdiblc2 = 1.044896747e-02 lpdiblc2 = -4.660380241e-9
+ pdiblcb = -0.025
+ drout = 3.009883541e-01 ldrout = 3.570453626e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.522960400e-07 lalpha0 = 5.885766851e-13 palpha0 = -1.323488980e-35
+ alpha1 = 0.85
+ beta0 = 1.208246472e+01 lbeta0 = 1.796707776e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.859191982e-01 lkt1 = -1.016563836e-8
+ kt2 = -2.530388930e-03 lkt2 = -2.418647259e-8
+ at = 2.628043600e+05 lat = -1.342367878e-1
+ ute = 6.275736411e-02 lute = -7.903188302e-7
+ ua1 = 4.049205174e-09 lua1 = -1.874859721e-15 pua1 = -8.271806126e-37
+ ub1 = -2.809220949e-18 lub1 = 1.461980805e-24
+ uc1 = -1.246391639e-11 luc1 = 6.067328922e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.168 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {2.303300179e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.774409178e-07 wvth0 = 1.155346505e-07 pvth0 = -5.901348198e-14
+ k1 = 2.296169368e-01 lk1 = 1.766711843e-07 wk1 = -4.134812492e-16 pk1 = 2.112003905e-22
+ k2 = -3.039964410e-02 lk2 = -7.365462557e-09 wk2 = 2.880021162e-08 pk2 = -1.471074489e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.763704446e+00 ldsub = -7.449717762e-07 wdsub = -5.048639779e-07 pdsub = 2.578774518e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446125e-03 lcdscd = -1.783892587e-09 wcdscd = -3.753421185e-18 pcdscd = 1.917195569e-24
+ cit = 0.0
+ voff = {-4.522962738e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.426031120e-07 wvoff = 8.883281999e-08 pvoff = -4.537456079e-14
+ nfactor = -8.485957432e+00 lnfactor = 5.194944330e-06 wnfactor = 3.233789858e-06 pnfactor = -1.651774586e-12
+ eta0 = 9.936117851e-01 leta0 = -2.572377985e-07 weta0 = 2.122630581e-09 peta0 = -1.084209984e-15
+ etab = 4.525776728e-02 letab = -2.327665454e-08 wetab = -1.785311287e-17 petab = 9.119109981e-24
+ u0 = 2.610173547e-02 lu0 = -3.265718191e-09 wu0 = -2.182443512e-09 pu0 = 1.114761592e-15
+ ua = -1.159362785e-09 lua = 2.013510626e-18 wua = -1.502971652e-17 pua = 7.676968781e-24
+ ub = 2.823582036e-18 lub = -8.794212960e-25 wub = -5.056896180e-25 pub = 2.582991772e-31
+ uc = -9.834907063e-11 luc = 5.248474075e-17 wuc = 3.366779216e-18 puc = -1.719703689e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.922456869e+04 lvsat = 1.410474085e-01 wvsat = 6.149494012e-02 pvsat = -3.141075449e-8
+ a0 = 1.500000004e+00 la0 = -2.288416567e-15 wa0 = -1.263108729e-15 pa0 = 6.451776891e-22
+ ags = -1.264024843e+00 lags = 6.556224824e-07 wags = -2.704426127e-16 pags = 1.381386082e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.842282574e-07 lb0 = 4.291257521e-13 wb0 = 2.151741894e-13 pb0 = -1.099079635e-19
+ b1 = -3.866595414e-07 lb1 = 2.041021896e-13 wb1 = 1.288488708e-13 pb1 = -6.581419934e-20
+ keta = 2.279719492e-01 lketa = -1.173389045e-07 wketa = -4.517171822e-08 pketa = 2.307308126e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.573701524e-01 lpclm = 8.366476370e-08 wpclm = 1.755862486e-07 ppclm = -8.968699758e-14
+ pdiblc1 = 6.485507005e-01 lpdiblc1 = -7.603960369e-08 wpdiblc1 = 2.162416912e-16 ppdiblc1 = -1.104530911e-22
+ pdiblc2 = -6.061561146e-03 lpdiblc2 = 3.772966630e-09 wpdiblc2 = -5.797922906e-18 ppdiblc2 = 2.961499102e-24
+ pdiblcb = 5.667376276e-02 lpdiblcb = -4.171781459e-08 wpdiblcb = -1.716726761e-17 ppdiblcb = 8.768791249e-24
+ drout = 1.518101819e+00 ldrout = -2.646391555e-07 wdrout = -1.145304296e-15 pdrout = 5.850055995e-22
+ pscbe1 = 8.089503011e+08 lpscbe1 = -4.571688497e+00 wpscbe1 = -1.131458282e-07 ppscbe1 = 5.779361725e-14
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.497450161e-06 lalpha0 = -4.584049782e-13 walpha0 = -9.173785118e-14 palpha0 = 4.685841005e-20
+ alpha1 = 0.85
+ beta0 = 1.771947945e+01 lbeta0 = -1.082600432e-06 wbeta0 = -2.446342721e-07 pbeta0 = 1.249557613e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.774161146e-01 lkt1 = -6.558749441e-08 wkt1 = -6.115856793e-08 pkt1 = 3.123894028e-14
+ kt2 = -7.179094734e-02 lkt2 = 1.119085100e-08 wkt2 = -6.862899138e-18 pkt2 = 3.505473689e-24
+ at = 1.170882334e+05 lat = -5.980703039e-02 wat = -4.586892592e-02 pat = 2.342920520e-8
+ ute = -1.264973424e+00 lute = -1.121325321e-07 wute = -1.223171357e-07 pute = 6.247788049e-14
+ ua1 = 7.985465814e-10 lua1 = -2.144688213e-16 wua1 = -1.294916094e-24 pua1 = 6.614250949e-31
+ ub1 = -6.300081721e-19 lub1 = 3.488694277e-25 wub1 = -1.839490838e-33 pub1 = 9.395863253e-40
+ uc1 = 6.369112720e-11 luc1 = 2.177435912e-17 wuc1 = 2.663459534e-26 puc1 = -1.360456199e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.169 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {1.981448708e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.792263209e-07 wvth0 = -4.126237517e-07 pvth0 = 7.872283510e-14
+ k1 = 9.070734848e-01 lk1 = 9.993081918e-16 wk1 = 1.476717415e-15 pk1 = -2.817370781e-22
+ k2 = 2.082612952e-01 lk2 = -6.960489427e-08 wk2 = -1.028578986e-07 pk2 = 1.962384705e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -5.771732862e+00 ldsub = 1.220164778e-06 wdsub = 1.803085635e-06 pdsub = -3.440034961e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999952e-03 lcdscd = 9.071346105e-18 wcdscd = 1.340508607e-17 pcdscd = -2.557501953e-24
+ cit = 0.0
+ voff = {9.177770648e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.146928337e-07 wvoff = -3.172600714e-07 pvoff = 6.052877998e-14
+ nfactor = 4.140333344e+01 lnfactor = -7.815484278e-06 wnfactor = -1.154924949e-05 pnfactor = 2.203435114e-12
+ eta0 = 2.688883937e-02 leta0 = -5.130013596e-09 weta0 = -7.580823504e-09 peta0 = 1.446314993e-15
+ etab = -4.399800023e-02 letab = 4.314765212e-17 wetab = 6.376105199e-17 petab = -1.216469980e-23
+ u0 = -6.646528651e-03 lu0 = 5.274570615e-09 wu0 = 7.794441116e-09 pu0 = -1.487070243e-15
+ ua = -1.290928864e-09 lua = 3.632410216e-17 wua = 5.367755899e-17 pua = -1.024092677e-23
+ ub = -5.235061817e-18 lub = 1.222160200e-24 wub = 1.806034350e-24 pub = -3.445660695e-31
+ uc = 1.341083321e-10 luc = -8.136895467e-18 wuc = -1.202421149e-17 puc = 2.294051213e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.031531142e+06 lvsat = -1.486221303e-01 wvsat = -2.196247862e-01 pvsat = 4.190133445e-8
+ a0 = 1.499999984e+00 la0 = 3.052702979e-15 wa0 = 4.511100826e-15 pa0 = -8.606546587e-22
+ ags = 1.249999997e+00 lags = 6.536122754e-16 wags = 9.658673861e-16 pags = -1.842739294e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.655394992e-06 lb0 = -5.200370366e-13 wb0 = -7.684792480e-13 pb0 = 1.466150818e-19
+ b1 = 1.590082190e-06 lb1 = -3.114043796e-13 wb1 = -4.601745387e-13 pb1 = 8.779485955e-20
+ keta = -6.405975466e-01 lketa = 1.091718600e-07 wketa = 1.613275651e-07 pketa = -3.077904083e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.405423034e+00 lpclm = -4.243601551e-07 wpclm = -6.270937450e-07 ppclm = 1.196407072e-13
+ pdiblc1 = 3.569721527e-01 lpdiblc1 = -5.226161726e-16 wpdiblc1 = -7.722906759e-16 ppdiblc1 = 1.473421385e-22
+ pdiblc2 = 8.406112027e-03 lpdiblc2 = 1.401253419e-17 wpdiblc2 = 2.070686678e-17 ppdiblc2 = -3.950582916e-24
+ pdiblcb = -1.032957702e-01 lpdiblcb = 4.149003363e-17 wpdiblcb = 6.131162245e-17 ppdiblcb = -1.169739305e-23
+ drout = 5.033266455e-01 ldrout = 2.767993390e-15 wdrout = 4.090373373e-15 pdrout = -7.803859781e-22
+ pscbe1 = 7.914198786e+08 lpscbe1 = 2.734546661e-07 wpscbe1 = 4.040946960e-07 ppscbe1 = -7.709574699e-14
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.110507114e-06 lalpha0 = 2.217137678e-13 walpha0 = 3.276351828e-13 palpha0 = -6.250820598e-20
+ alpha1 = 0.85
+ beta0 = 1.130104767e+01 lbeta0 = 5.912367196e-07 wbeta0 = 8.736938288e-07 pbeta0 = -1.666885508e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.956988219e-01 lkt1 = 1.478091797e-07 wkt1 = 2.184234569e-07 pkt1 = -4.167213765e-14
+ kt2 = -2.887893909e-02 lkt2 = 1.658642668e-17 wkt2 = 2.451039371e-17 pkt2 = -4.676245502e-24
+ at = -5.373330741e+05 lat = 1.108568847e-01 wat = 1.638175926e-01 pat = -3.125410322e-8
+ ute = -2.828519362e+00 lute = 2.956183591e-07 wute = 4.368469133e-07 pute = -8.334427521e-14
+ ua1 = -2.384735240e-11 lua1 = 3.129577774e-24 wua1 = 4.624700579e-24 pua1 = -8.823281236e-31
+ ub1 = 7.077531467e-19 lub1 = 4.445715765e-33 wub1 = 6.569610508e-33 pub1 = -1.253389623e-39
+ uc1 = 1.471862503e-10 luc1 = -6.437098847e-26 wuc1 = -9.512349570e-26 puc1 = 1.814823924e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.170 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {-1.307351324e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.237487853e-07 wvth0 = 1.795588670e-07 pvth0 = -3.425731800e-14
+ k1 = 0.90707349
+ k2 = 9.806228507e-02 lk2 = -4.858046592e-08 wk2 = -6.719062103e-08 pk2 = 1.281902982e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.429490745e+00 ldsub = -5.352998694e-07 wdsub = -8.752065606e-07 pdsub = 1.669771589e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = -1.343760374e+01 lnfactor = 2.647398761e-06 wnfactor = 1.621325400e-06 pnfactor = -3.093261878e-13
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = 1.766145641e-01 lu0 = -2.968908023e-08 wu0 = -6.587716269e-08 pu0 = 1.256844036e-14
+ ua = -1.072899214e-09 lua = -5.272902601e-18 wua = 1.329021165e-16 pua = -2.535586320e-23
+ ub = -6.163090404e-18 lub = 1.399215062e-24 wub = 5.016658097e-25 pub = -9.571081316e-32
+ uc = -1.113153575e-10 luc = 3.868650857e-17 wuc = 1.020478326e-16 puc = -1.946929779e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.306845638e+05 lvsat = 7.311235533e-02 wvsat = 1.016641890e-01 pvsat = -1.939610396e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.055917419e-06 lb0 = -5.964511084e-13 wb0 = -3.644689769e-13 pb0 = 6.953557823e-20
+ b1 = 2.309490899e-06 lb1 = -4.486574896e-13 wb1 = -1.372673939e-12 pb1 = 2.618869702e-19
+ keta = -1.131181136e+00 lketa = 2.027683406e-07 wketa = 3.716864939e-07 pketa = -7.091257942e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.438503395e-02 lpclm = 2.990856081e-08 wpclm = 1.113922654e-07 ppclm = -2.125208474e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.673659118e-07 lalpha0 = -2.208651526e-14 walpha0 = 2.542867870e-21 palpha0 = -4.851435998e-28
+ alpha1 = 0.85
+ beta0 = 1.734774328e+01 lbeta0 = -5.623881488e-07 wbeta0 = 1.759190127e-14 pbeta0 = -3.356277034e-21
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.137700705e-01 lkt1 = -2.045047907e-08 wkt1 = -8.760734360e-16 pkt1 = 1.671425220e-22
+ kt2 = -0.028878939
+ at = -9.874845431e+03 lat = 1.022523909e-02 wat = -2.813644242e-10 pat = 5.368038546e-17
+ ute = -9.888383039e-01 lute = -5.536703130e-08 wute = -1.908327907e-07 pute = 3.640822481e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.171 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.481164+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.031936246
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.9222
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0220043
+ ua = -1.0491453e-9
+ ub = 1.24835e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.4304e-8
+ b1 = 1.2375e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.172 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.627150263e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.691784641e-7
+ k1 = 5.566262089e-01 lk1 = 2.277529835e-7
+ k2 = -2.165726269e-02 lk2 = -2.056905354e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017327274e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.309728469e-7
+ nfactor = 4.223472310e+00 lnfactor = -6.028695726e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.069834161e-02 lu0 = 2.613325382e-8
+ ua = -1.131262846e-09 lua = 1.643236638e-15
+ ub = 1.288370552e-18 lub = -8.008426962e-25
+ uc = 6.338098646e-11 luc = -2.970398364e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.479156936e+00 la0 = -2.332395909e-6
+ ags = 3.213416405e-01 lags = 4.710210753e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.387376907e-08 lb0 = 1.914986009e-13
+ b1 = 1.774850174e-08 lb1 = -1.075279933e-13
+ keta = -1.957380452e-03 lketa = -5.181231829e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.762224597e-02 lpclm = 8.904248667e-07 ppclm = -1.110223025e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.597527482e-04 lpdiblc2 = 2.241368535e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -6.737507727e+07 lpscbe1 = 5.850655103e+03 ppscbe1 = -9.536743164e-19
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.784760245e-01 lkt1 = -1.581647627e-7
+ kt2 = -2.846385108e-02 lkt2 = -2.109296763e-8
+ at = 1.883513100e+05 lat = -2.671702072e-1
+ ute = -1.123944838e+00 lute = 1.709889326e-7
+ ua1 = 8.756696787e-10 lua1 = 4.909252558e-15
+ ub1 = -2.470825931e-19 lub1 = -6.451225409e-24
+ uc1 = 4.320065665e-11 luc1 = -1.877470904e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.173 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {4.960531199e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.021141305e-7
+ k1 = 6.074825579e-01 lk1 = -1.796463452e-7
+ k2 = -5.290211314e-02 lk2 = 4.460527524e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.260637441e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.393772087e-8
+ nfactor = 4.057176644e+00 lnfactor = -4.696536728e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.133884946e-02 lu0 = 2.100228251e-8
+ ua = -1.247236071e-09 lua = 2.572273326e-15
+ ub = 1.471300791e-18 lub = -2.266257692e-24
+ uc = 3.261899065e-11 luc = -5.061207102e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.206048537e+00 la0 = -1.445829675e-7
+ ags = 4.068117269e-01 lags = -2.136614964e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.372805585e-08 lb0 = -4.301530117e-13 wb0 = -8.530300067e-31 pb0 = 2.874452629e-35
+ b1 = 3.316787051e-09 lb1 = 8.081384646e-15
+ keta = -1.933584143e-02 lketa = 8.740281358e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.490412944e-01 lpclm = 3.465244080e-06 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.079775722e-03 lpdiblc2 = 2.978379250e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.255747443e+08 lpscbe1 = 1.100660974e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.825979885e-01 lkt1 = -1.251445908e-7
+ kt2 = -1.846134680e-02 lkt2 = -1.012208889e-7
+ at = 1.700404475e+05 lat = -1.204858063e-1
+ ute = -8.041975216e-01 lute = -2.390438396e-6
+ ua1 = 2.400933761e-09 lua1 = -7.309311599e-15
+ ub1 = -1.693975356e-18 lub1 = 5.139522876e-24
+ uc1 = -1.227453723e-11 luc1 = 2.566528161e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.174 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.099735415e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.628229852e-8
+ k1 = 5.212762443e-01 lk1 = 1.661087306e-7
+ k2 = -2.315691021e-02 lk2 = -7.469636824e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.116123628e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.976323031e-9
+ nfactor = 2.892332897e+00 lnfactor = -2.459773863e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.846443345e-02 lu0 = -7.576909981e-9
+ ua = -4.928630170e-10 lua = -4.533555576e-16
+ ub = 8.765807986e-19 lub = 1.190369253e-25
+ uc = -5.592278815e-12 luc = 1.026451536e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.163327600e+04 lvsat = 2.742042995e-1
+ a0 = 8.382203100e-01 la0 = 1.330697336e-6
+ ags = 4.391592679e-01 lags = -3.434005609e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.133074850e-10 lb0 = -2.163189654e-13
+ b1 = -3.280798056e-09 lb1 = 3.454288663e-14
+ keta = -1.309633638e-02 lketa = 6.237749411e-08 wketa = 1.734723476e-24
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.744363068e-01 lpclm = 5.171412440e-06 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -7.611070267e-04 lpdiblc2 = 2.850568056e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.055457235e-01 lkt1 = -3.310613675e-8
+ kt2 = -5.702681193e-02 lkt2 = 5.345693870e-08 wkt2 = -2.775557562e-23
+ at = 140000.0
+ ute = -1.616761652e+00 lute = 8.685824428e-7
+ ua1 = -3.410928692e-10 lua1 = 3.688370421e-15
+ ub1 = 6.948567385e-20 lub1 = -1.933341932e-24
+ uc1 = 5.824216620e-11 luc1 = -2.617459078e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.175 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.069953072e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.227089047e-8
+ k1 = 6.223438819e-01 lk1 = -3.711666019e-8
+ k2 = -6.443184982e-02 lk2 = 8.298702475e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.632358000e-01 ldsub = -6.097423013e-07 wdsub = -4.440892099e-22
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.759591720e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.220774955e-8
+ nfactor = 3.211669446e+00 lnfactor = -6.667151992e-7
+ eta0 = 1.583043279e-01 leta0 = -1.574532464e-7
+ etab = -1.404391494e-01 letab = 1.416380554e-7
+ u0 = 2.973415850e-02 lu0 = -1.013005535e-08 wu0 = -1.387778781e-23
+ ua = -2.241512811e-10 lua = -9.936773541e-16
+ ub = 5.476179603e-19 lub = 7.805107952e-25
+ uc = 4.840043040e-11 luc = -5.922630220e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.196979920e+05 lvsat = 5.690928146e-2
+ a0 = 1.5
+ ags = 3.352030625e-01 lags = -1.343668785e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.321102943e-07 lb0 = -4.811334227e-13 pb0 = -1.058791184e-34
+ b1 = 5.641899952e-09 lb1 = 1.660125039e-14
+ keta = 1.805777867e-02 lketa = -2.667642893e-10
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.567618932e+00 lpclm = -1.548745445e-6
+ pdiblc1 = 1.884437022e-01 lpdiblc1 = 4.052865819e-7
+ pdiblc2 = 2.107396742e-02 lpdiblc2 = -1.539998143e-8
+ pdiblcb = -0.025
+ drout = 4.647599830e-01 ldrout = 1.915072929e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.483244388e-01 lkt1 = 5.291270522e-8
+ kt2 = -3.446762206e-02 lkt2 = 8.095235534e-9
+ at = 1.501078600e+05 lat = -2.032474338e-2
+ ute = -1.655494688e+00 lute = 9.464662882e-7
+ ua1 = 7.844854756e-10 lua1 = 1.425073244e-15
+ ub1 = -4.160807111e-19 lub1 = -9.569718432e-25
+ uc1 = 4.286300461e-11 luc1 = 4.749612046e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.176 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {5.392887653e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.962911505e-8
+ k1 = 5.959670436e-01 lk1 = -1.045532135e-8
+ k2 = -6.786986822e-02 lk2 = 1.177380334e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.138011941e-01 ldsub = 4.669710627e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.486568763e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.529100738e-8
+ nfactor = 3.438318471e+00 lnfactor = -8.958088615e-7
+ eta0 = -4.954531759e-01 leta0 = 5.033556859e-07 weta0 = -1.214306433e-23 peta0 = -7.112366252e-29
+ etab = -0.0003125
+ u0 = 1.971626586e-02 lu0 = -4.109710889e-12
+ ua = -1.260147125e-09 lua = 5.349274039e-17
+ ub = 1.542420970e-18 lub = -2.250221600e-25
+ uc = 8.150086973e-11 luc = -3.938009089e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.546354561e+05 lvsat = 2.159498183e-2
+ a0 = 1.5
+ ags = 3.889507903e-01 lags = -1.886943293e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.479878483e-07 lb0 = 2.063002585e-13
+ b1 = 3.140418965e-08 lb1 = -9.438911366e-15
+ keta = 3.775962016e-02 lketa = -2.018110984e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.458569580e+00 lpclm = -4.277338871e-7
+ pdiblc1 = 6.810636468e-01 lpdiblc1 = -9.264676145e-8
+ pdiblc2 = 1.044896747e-02 lpdiblc2 = -4.660380241e-9
+ pdiblcb = -0.025
+ drout = 3.009883541e-01 ldrout = 3.570453626e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.522960400e-07 lalpha0 = 5.885766851e-13 walpha0 = -5.293955920e-29 palpha0 = 1.058791184e-34
+ alpha1 = 0.85
+ beta0 = 1.208246472e+01 lbeta0 = 1.796707776e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.859191982e-01 lkt1 = -1.016563836e-8
+ kt2 = -2.530388930e-03 lkt2 = -2.418647259e-8
+ at = 2.628043600e+05 lat = -1.342367878e-1
+ ute = 6.275736411e-02 lute = -7.903188302e-7
+ ua1 = 4.049205174e-09 lua1 = -1.874859721e-15
+ ub1 = -2.809220949e-18 lub1 = 1.461980805e-24
+ uc1 = -1.246391639e-11 luc1 = 6.067328922e-17 puc1 = 1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.177 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {6.401261761e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.187722263e-8
+ k1 = 2.296169353e-01 lk1 = 1.766711851e-7
+ k2 = 7.175339854e-02 lk2 = -5.954380660e-08 pk2 = 6.938893904e-30
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -2.702515522e-02 ldsub = 1.697078339e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.892446112e-03 lcdscd = -1.783892580e-9
+ cit = 0.0
+ voff = {-1.372102957e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.833839441e-8
+ nfactor = 2.984148331e+00 lnfactor = -6.638251119e-7
+ eta0 = 1.001140660e+00 leta0 = -2.610834421e-7
+ etab = 4.525776721e-02 letab = -2.327665451e-08 wetab = 1.517883041e-24 petab = -2.602085214e-30
+ u0 = 1.836070744e-02 lu0 = 6.882905486e-10
+ ua = -1.212672507e-09 lua = 2.924337024e-17
+ ub = 1.029923927e-18 lub = 3.675415476e-26
+ uc = -8.640725765e-11 luc = 4.638502987e-17 wuc = 6.462348536e-33 puc = 8.077935669e-40
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.388951911e+05 lvsat = 2.963488884e-2
+ a0 = 1.5
+ ags = -1.264024844e+00 lags = 6.556224829e-07 wags = -2.081668171e-22 pags = -5.898059818e-29
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.210151797e-07 lb0 = 3.928719698e-14 wb0 = 1.058791184e-28
+ b1 = 7.036155178e-08 lb1 = -2.933778654e-14 wb1 = -1.323488980e-29 pb1 = -6.617444900e-36
+ keta = 6.774991616e-02 lketa = -3.549973317e-08 wketa = -1.387778781e-23 pketa = -2.602085214e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.080166602e+00 lpclm = -2.344509436e-7
+ pdiblc1 = 6.485507013e-01 lpdiblc1 = -7.603960408e-8
+ pdiblc2 = -6.061561167e-03 lpdiblc2 = 3.772966640e-09 ppdiblc2 = 2.168404345e-31
+ pdiblcb = 5.667376270e-02 lpdiblcb = -4.171781455e-8
+ drout = 1.518101815e+00 ldrout = -2.646391535e-7
+ pscbe1 = 8.089503007e+08 lpscbe1 = -4.571688292e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.172060170e-06 lalpha0 = -2.922003258e-13
+ alpha1 = 0.85
+ beta0 = 1.685177280e+01 lbeta0 = -6.393880214e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.943427775e-01 lkt1 = 4.521560804e-8
+ kt2 = -7.179094737e-02 lkt2 = 1.119085101e-8
+ at = -4.560676369e+04 lat = 2.329529640e-2
+ ute = -1.698826749e+00 lute = 1.094736726e-7
+ ua1 = 7.985465768e-10 lua1 = -2.144688189e-16 wua1 = -2.067951531e-31
+ ub1 = -6.300081786e-19 lub1 = 3.488694311e-25 wub1 = 9.629649722e-41 pub1 = -1.203706215e-47
+ uc1 = 6.369112730e-11 luc1 = 2.177435907e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.178 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {0.517891+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = -0.156571
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.62373
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 0.43867
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = 0.021
+ ua = -1.100537e-9
+ ub = 1.17086e-18
+ uc = 9.1459e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 252532.0
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.0366e-8
+ b1 = -4.2136e-8
+ keta = -0.068376
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.18115
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.16e-8
+ alpha1 = 0.85
+ beta0 = 14.4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.22096074
+ kt2 = -0.028878939
+ at = 43720.487
+ ute = -1.2790432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.179 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.363696e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.052*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 5.4034e-8
+ lint = -5.393e-9
+ vth0 = {-5.540233200e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.045062455e-07 wvth0 = 2.988973523e-07 pvth0 = -5.702543026e-14
+ k1 = 0.90707349
+ k2 = -2.325260563e-01 lk2 = 1.449116137e-08 wk2 = 2.601281122e-08 pk2 = -4.962880202e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.308003241e+00 ldsub = -5.121217546e-07 wdsub = -8.409553457e-07 pdsub = 1.604425066e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = -1.343760560e+01 lnfactor = 2.647399117e-06 wnfactor = 1.621325926e-06 pnfactor = -3.093262881e-13
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = -1.159522987e-02 lu0 = 6.218713526e-09 wu0 = -1.281479905e-08 pu0 = 2.444884252e-15
+ ua = -1.072897415e-09 lua = -5.273245830e-18 wua = 1.329016093e-16 pua = -2.535576643e-23
+ ub = -6.163134324e-18 lub = 1.399223441e-24 wub = 5.016781923e-25 pub = -9.571317560e-32
+ uc = -9.715009267e-11 luc = 3.598397435e-17 wuc = 9.805419118e-17 puc = -1.870736692e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.616972904e+05 lvsat = -7.806300910e-02 wvsat = -1.217336119e-01 pvsat = 2.322506889e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.055925333e-06 lb0 = -5.964526183e-13 wb0 = -3.644712082e-13 pb0 = 6.953600393e-20
+ b1 = 2.309501807e-06 lb1 = -4.486595707e-13 wb1 = -1.372677015e-12 pb1 = 2.618875569e-19
+ keta = -1.131181040e+00 lketa = 2.027683223e-07 wketa = 3.716864668e-07 pketa = -7.091257426e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.438497216e-02 lpclm = 2.990857260e-08 wpclm = 1.113922828e-07 ppclm = -2.125208807e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.673659202e-07 lalpha0 = -2.208651686e-14 walpha0 = 1.811849002e-22 palpha0 = -3.456754693e-29
+ alpha1 = 0.85
+ beta0 = 1.734774334e+01 lbeta0 = -5.623881607e-07 wbeta0 = 3.171862772e-17 pbeta0 = -6.053824109e-24
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -6.928e-9
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 2.4384e-10
+ cgdo = 2.4384e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00163782571
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 4.49076474e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.91230478e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.137700734e-01 lkt1 = -2.045047852e-08 wkt1 = -6.743006153e-17 pkt1 = 1.286470930e-23
+ kt2 = -0.028878939
+ at = -9.874846353e+03 lat = 1.022523927e-02 wat = -2.139387652e-11 pat = 4.081666702e-18
+ ute = -1.015327828e+00 lute = -5.031320101e-08 wute = -1.833645463e-07 pute = 3.498338833e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
.ends sky130_fd_pr__nfet_01v8
* Well Proximity Effect Parameters
